##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Tue Oct 27 22:00:12 2020
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO temp_wrapper
  CLASS BLOCK ;
  SIZE 2078.280000 BY 2078.080000 ;
  FOREIGN temp_wrapper 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN RESET_REGn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.7884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 17.766 LAYER met3  ;
    ANTENNAMAXAREACAR 10.4844 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.6182 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.125802 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 384.642 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2054.24 LAYER met4  ;
    ANTENNAGATEAREA 947.52 LAYER met4  ;
    ANTENNAMAXAREACAR 32.4314 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 161.604 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.500997 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 189.180000 0.800000 189.480000 ;
    END
  END RESET_REGn
  PIN SEL_CONV_TIME_REG[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 336.405 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1798.37 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 9.423 LAYER met3  ;
    ANTENNAMAXAREACAR 112.51 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 571.006 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.412489 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 234.184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1251.33 LAYER met4  ;
    ANTENNAGATEAREA 33.696 LAYER met4  ;
    ANTENNAMAXAREACAR 120.191 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 611.581 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.435559 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 378.280000 0.800000 378.580000 ;
    END
  END SEL_CONV_TIME_REG[3]
  PIN SEL_CONV_TIME_REG[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1033.57 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5530.18 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 56.889 LAYER met3  ;
    ANTENNAMAXAREACAR 70.1185 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 351.733 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.542416 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 80.4975 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 430.256 LAYER met4  ;
    ANTENNAGATEAREA 77.472 LAYER met4  ;
    ANTENNAMAXAREACAR 71.1575 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 358.735 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.542416 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 566.770000 0.800000 567.070000 ;
    END
  END SEL_CONV_TIME_REG[2]
  PIN SEL_CONV_TIME_REG[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 359.376 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1922.26 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 48.672 LAYER met3  ;
    ANTENNAMAXAREACAR 79.2607 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 395.615 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.461846 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 90.3372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 478.584 LAYER met4  ;
    ANTENNAGATEAREA 86.022 LAYER met4  ;
    ANTENNAMAXAREACAR 80.3109 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 401.179 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.469286 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 116.272 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 178.248 LAYER met5  ;
    ANTENNAGATEAREA 113.184 LAYER met5  ;
    ANTENNAMAXAREACAR 81.3381 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 424.821 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 755.870000 0.800000 756.170000 ;
    END
  END SEL_CONV_TIME_REG[1]
  PIN SEL_CONV_TIME_REG[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 797.629 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4263.37 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 53.928 LAYER met3  ;
    ANTENNAMAXAREACAR 53.5513 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 269.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.375514 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 153.476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 819.472 LAYER met4  ;
    ANTENNAGATEAREA 88.416 LAYER met4  ;
    ANTENNAMAXAREACAR 55.2871 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 278.517 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.426692 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 944.360000 0.800000 944.660000 ;
    END
  END SEL_CONV_TIME_REG[0]
  PIN CLK_REF
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 184.311 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 983.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.576 LAYER met4  ;
    ANTENNAMAXAREACAR 4.69358 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 24.9583 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.228125 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 0.690000 0.800000 0.990000 ;
    END
  END CLK_REF
  PIN SEL_DESIGN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.052 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.88 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.305 LAYER met3  ;
    ANTENNAMAXAREACAR 52.4669 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 268.231 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1133.460000 0.800000 1133.760000 ;
    END
  END SEL_DESIGN
  PIN SEL_GROUP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.3424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8 LAYER met3  ;
    ANTENNAMAXAREACAR 65.4575 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 326.368 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.229899 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1321.950000 0.800000 1322.250000 ;
    END
  END SEL_GROUP[2]
  PIN SEL_GROUP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.291 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8 LAYER met3  ;
    ANTENNAMAXAREACAR 12.5856 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 60.1353 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.530909 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1511.050000 0.800000 1511.350000 ;
    END
  END SEL_GROUP[1]
  PIN SEL_GROUP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.176 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0475 LAYER met3  ;
    ANTENNAMAXAREACAR 50.5838 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 252.106 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.278788 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1699.540000 0.800000 1699.840000 ;
    END
  END SEL_GROUP[0]
  PIN SEL_INST[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.6566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 186.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0575 LAYER met3  ;
    ANTENNAMAXAREACAR 34.596 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 183.187 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1888.640000 0.800000 1888.940000 ;
    END
  END SEL_INST[1]
  PIN SEL_INST[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.3738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 180.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.485 LAYER met3  ;
    ANTENNAMAXAREACAR 24.5636 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.752 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2077.740000 0.800000 2078.040000 ;
    END
  END SEL_INST[0]
  PIN CLK_OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.9504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1994.780000 2078.280000 1995.080000 ;
    END
  END CLK_OUT
  PIN DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.6344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 232.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1911.820000 2078.280000 1912.120000 ;
    END
  END DOUT[23]
  PIN DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1828.860000 2078.280000 1829.160000 ;
    END
  END DOUT[22]
  PIN DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.7004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.064 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1745.900000 2078.280000 1746.200000 ;
    END
  END DOUT[21]
  PIN DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.1214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1662.330000 2078.280000 1662.630000 ;
    END
  END DOUT[20]
  PIN DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 49.6392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 265.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1579.370000 2078.280000 1579.670000 ;
    END
  END DOUT[19]
  PIN DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 53.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 285.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1496.410000 2078.280000 1496.710000 ;
    END
  END DOUT[18]
  PIN DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.0324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1413.450000 2078.280000 1413.750000 ;
    END
  END DOUT[17]
  PIN DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.3634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1330.490000 2078.280000 1330.790000 ;
    END
  END DOUT[16]
  PIN DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.3314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 199.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1246.920000 2078.280000 1247.220000 ;
    END
  END DOUT[15]
  PIN DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 52.0332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1163.960000 2078.280000 1164.260000 ;
    END
  END DOUT[14]
  PIN DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 114.73 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 612.36 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1081.000000 2078.280000 1081.300000 ;
    END
  END DOUT[13]
  PIN DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 42.3924 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 998.040000 2078.280000 998.340000 ;
    END
  END DOUT[12]
  PIN DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.8584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.24 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 915.080000 2078.280000 915.380000 ;
    END
  END DOUT[11]
  PIN DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 142.975 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 763 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 831.510000 2078.280000 831.810000 ;
    END
  END DOUT[10]
  PIN DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 230.216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1227.81 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.096 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.7155 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 205.264 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 311.736 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 748.550000 2078.280000 748.850000 ;
    END
  END DOUT[9]
  PIN DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 269.65 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1438.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 665.590000 2078.280000 665.890000 ;
    END
  END DOUT[8]
  PIN DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.2194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 107.832 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 582.630000 2078.280000 582.930000 ;
    END
  END DOUT[7]
  PIN DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.4964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 499.670000 2078.280000 499.970000 ;
    END
  END DOUT[6]
  PIN DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7155 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.8114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 416.710000 2078.280000 417.010000 ;
    END
  END DOUT[5]
  PIN DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.3634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 333.140000 2078.280000 333.440000 ;
    END
  END DOUT[4]
  PIN DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.7324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 250.180000 2078.280000 250.480000 ;
    END
  END DOUT[3]
  PIN DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7952 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.4674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 178.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 167.220000 2078.280000 167.520000 ;
    END
  END DOUT[2]
  PIN DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.9424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 84.260000 2078.280000 84.560000 ;
    END
  END DOUT[1]
  PIN DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.128 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 1.300000 2078.280000 1.600000 ;
    END
  END DOUT[0]
  PIN DONE
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.4674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 178.488 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2077.480000 2077.740000 2078.280000 2078.040000 ;
    END
  END DONE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2044.780000 2066.880000 2055.980000 2078.080000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.780000 0.000000 2055.980000 11.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 22.300000 2066.880000 33.500000 2078.080000 ;
    END
    PORT
      LAYER met4 ;
        RECT 22.300000 0.000000 33.500000 11.200000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2067.080000 2043.900000 2078.280000 2055.100000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2043.900000 11.200000 2055.100000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2067.080000 22.300000 2078.280000 33.500000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 22.300000 11.200000 33.500000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 1039.100000 39.100000 1042.300000 2038.300000 ;
        RECT 22.300000 0.000000 33.500000 2078.080000 ;
        RECT 274.100000 39.100000 277.300000 2038.300000 ;
        RECT 499.100000 39.100000 502.300000 2038.300000 ;
        RECT 539.100000 39.100000 542.300000 2038.300000 ;
        RECT 774.100000 39.100000 777.300000 2038.300000 ;
        RECT 1009.100000 39.100000 1012.300000 2038.300000 ;
        RECT 146.940000 1019.100000 148.540000 1090.640000 ;
        RECT 241.500000 1019.100000 243.100000 1090.640000 ;
        RECT 338.780000 1019.100000 340.380000 1090.640000 ;
        RECT 439.580000 1019.100000 441.180000 1090.640000 ;
        RECT 636.860000 1019.100000 638.460000 1090.640000 ;
        RECT 731.420000 1019.100000 733.020000 1090.640000 ;
        RECT 828.700000 1019.100000 830.300000 1090.640000 ;
        RECT 929.500000 1019.100000 931.100000 1090.640000 ;
        RECT 2044.780000 0.000000 2055.980000 2078.080000 ;
        RECT 1274.100000 39.100000 1277.300000 2038.300000 ;
        RECT 1519.100000 39.100000 1522.300000 2038.300000 ;
        RECT 1539.100000 39.100000 1542.300000 2038.300000 ;
        RECT 1774.100000 39.100000 1777.300000 2038.300000 ;
        RECT 2029.100000 39.100000 2032.300000 2038.300000 ;
        RECT 1622.940000 1019.100000 1624.540000 1090.640000 ;
        RECT 1717.500000 1019.100000 1719.100000 1090.640000 ;
        RECT 1814.780000 1019.100000 1816.380000 1090.640000 ;
        RECT 1915.580000 1019.100000 1917.180000 1090.640000 ;
        RECT 1126.780000 1019.100000 1128.380000 1096.560000 ;
        RECT 1227.580000 1019.100000 1229.180000 1096.560000 ;
        RECT 1324.860000 1019.100000 1326.460000 1096.560000 ;
        RECT 1425.660000 1019.100000 1427.260000 1096.560000 ;
        RECT 1039.100000 22.300000 1042.300000 39.100000 ;
        RECT 241.500000 250.410000 243.100000 282.300000 ;
        RECT 439.580000 256.330000 441.180000 282.300000 ;
        RECT 241.500000 22.300000 243.100000 139.900000 ;
        RECT 146.940000 22.300000 148.540000 139.900000 ;
        RECT 439.580000 22.300000 441.180000 139.900000 ;
        RECT 338.780000 22.300000 340.380000 139.900000 ;
        RECT 274.100000 22.300000 277.300000 39.100000 ;
        RECT 499.100000 22.300000 502.300000 39.100000 ;
        RECT 247.740000 279.100000 249.340000 332.010000 ;
        RECT 146.940000 279.100000 148.540000 332.010000 ;
        RECT 247.740000 448.440000 249.340000 472.300000 ;
        RECT 146.940000 448.440000 148.540000 472.300000 ;
        RECT 338.780000 279.100000 340.380000 332.010000 ;
        RECT 439.580000 279.100000 441.180000 332.010000 ;
        RECT 439.580000 448.440000 441.180000 472.300000 ;
        RECT 731.420000 250.410000 733.020000 282.300000 ;
        RECT 929.500000 256.330000 931.100000 282.300000 ;
        RECT 828.700000 256.330000 830.300000 282.300000 ;
        RECT 731.420000 22.300000 733.020000 139.900000 ;
        RECT 636.860000 22.300000 638.460000 139.900000 ;
        RECT 539.100000 22.300000 542.300000 39.100000 ;
        RECT 774.100000 22.300000 777.300000 39.100000 ;
        RECT 929.500000 22.300000 931.100000 139.900000 ;
        RECT 828.700000 22.300000 830.300000 139.900000 ;
        RECT 1009.100000 22.300000 1012.300000 39.100000 ;
        RECT 636.860000 279.100000 638.460000 332.010000 ;
        RECT 737.660000 279.100000 739.260000 332.010000 ;
        RECT 737.660000 448.440000 739.260000 472.300000 ;
        RECT 828.700000 279.100000 830.300000 332.010000 ;
        RECT 929.500000 279.100000 931.100000 332.010000 ;
        RECT 828.700000 448.440000 830.300000 472.300000 ;
        RECT 929.500000 448.440000 931.100000 472.300000 ;
        RECT 421.780000 769.100000 423.380000 810.340000 ;
        RECT 338.780000 769.100000 340.380000 810.340000 ;
        RECT 229.940000 769.100000 231.540000 810.340000 ;
        RECT 146.940000 769.100000 148.540000 810.340000 ;
        RECT 229.940000 529.100000 231.540000 630.040000 ;
        RECT 146.940000 529.100000 148.540000 630.040000 ;
        RECT 229.940000 728.740000 231.540000 772.300000 ;
        RECT 338.780000 529.100000 340.380000 630.040000 ;
        RECT 421.780000 529.100000 423.380000 630.040000 ;
        RECT 338.780000 728.740000 340.380000 772.300000 ;
        RECT 421.780000 728.740000 423.380000 772.300000 ;
        RECT 229.940000 909.040000 231.540000 952.300000 ;
        RECT 146.940000 909.040000 148.540000 952.300000 ;
        RECT 421.780000 909.040000 423.380000 952.300000 ;
        RECT 338.780000 909.040000 340.380000 952.300000 ;
        RECT 911.700000 769.100000 913.300000 810.340000 ;
        RECT 828.700000 769.100000 830.300000 810.340000 ;
        RECT 719.860000 769.100000 721.460000 810.340000 ;
        RECT 636.860000 769.100000 638.460000 810.340000 ;
        RECT 636.860000 529.100000 638.460000 630.040000 ;
        RECT 719.860000 529.100000 721.460000 630.040000 ;
        RECT 719.860000 728.740000 721.460000 772.300000 ;
        RECT 828.700000 529.100000 830.300000 630.040000 ;
        RECT 911.700000 529.100000 913.300000 630.040000 ;
        RECT 828.700000 728.740000 830.300000 772.300000 ;
        RECT 911.700000 728.740000 913.300000 772.300000 ;
        RECT 719.860000 909.040000 721.460000 952.300000 ;
        RECT 828.700000 909.040000 830.300000 952.300000 ;
        RECT 911.700000 909.040000 913.300000 952.300000 ;
        RECT 1425.660000 256.330000 1427.260000 282.300000 ;
        RECT 1324.860000 256.330000 1326.460000 282.300000 ;
        RECT 1227.580000 256.330000 1229.180000 282.300000 ;
        RECT 1227.580000 22.300000 1229.180000 139.900000 ;
        RECT 1126.780000 22.300000 1128.380000 139.900000 ;
        RECT 1274.100000 22.300000 1277.300000 39.100000 ;
        RECT 1425.660000 22.300000 1427.260000 139.900000 ;
        RECT 1324.860000 22.300000 1326.460000 139.900000 ;
        RECT 1519.100000 22.300000 1522.300000 39.100000 ;
        RECT 1539.100000 22.300000 1542.300000 39.100000 ;
        RECT 1126.780000 279.100000 1128.380000 337.930000 ;
        RECT 1227.580000 279.100000 1229.180000 337.930000 ;
        RECT 1126.780000 454.360000 1128.380000 472.300000 ;
        RECT 1227.580000 454.360000 1229.180000 472.300000 ;
        RECT 1425.660000 279.100000 1427.260000 337.930000 ;
        RECT 1324.860000 279.100000 1326.460000 337.930000 ;
        RECT 1425.660000 454.360000 1427.260000 472.300000 ;
        RECT 1324.860000 454.360000 1326.460000 472.300000 ;
        RECT 1717.500000 250.410000 1719.100000 282.300000 ;
        RECT 1915.580000 256.330000 1917.180000 282.300000 ;
        RECT 1814.780000 256.330000 1816.380000 282.300000 ;
        RECT 1814.780000 22.300000 1816.380000 139.900000 ;
        RECT 1717.500000 22.300000 1719.100000 139.900000 ;
        RECT 1622.940000 22.300000 1624.540000 139.900000 ;
        RECT 1774.100000 22.300000 1777.300000 39.100000 ;
        RECT 1915.580000 22.300000 1917.180000 139.900000 ;
        RECT 2029.100000 22.300000 2032.300000 39.100000 ;
        RECT 1622.940000 279.100000 1624.540000 332.010000 ;
        RECT 1723.740000 279.100000 1725.340000 332.010000 ;
        RECT 1814.780000 279.100000 1816.380000 332.010000 ;
        RECT 1814.780000 448.440000 1816.380000 472.300000 ;
        RECT 1723.740000 448.440000 1725.340000 472.300000 ;
        RECT 1915.580000 279.100000 1917.180000 332.010000 ;
        RECT 1915.580000 448.440000 1917.180000 472.300000 ;
        RECT 1407.860000 769.100000 1409.460000 816.260000 ;
        RECT 1324.860000 769.100000 1326.460000 816.260000 ;
        RECT 1209.780000 769.100000 1211.380000 816.260000 ;
        RECT 1126.780000 769.100000 1128.380000 816.260000 ;
        RECT 1126.780000 529.100000 1128.380000 635.960000 ;
        RECT 1209.780000 529.100000 1211.380000 635.960000 ;
        RECT 1209.780000 734.660000 1211.380000 772.300000 ;
        RECT 1407.860000 529.100000 1409.460000 635.960000 ;
        RECT 1324.860000 529.100000 1326.460000 635.960000 ;
        RECT 1324.860000 734.660000 1326.460000 772.300000 ;
        RECT 1407.860000 734.660000 1409.460000 772.300000 ;
        RECT 1126.780000 914.960000 1128.380000 952.300000 ;
        RECT 1209.780000 914.960000 1211.380000 952.300000 ;
        RECT 1324.860000 914.960000 1326.460000 952.300000 ;
        RECT 1407.860000 914.960000 1409.460000 952.300000 ;
        RECT 1897.780000 769.100000 1899.380000 810.340000 ;
        RECT 1814.780000 769.100000 1816.380000 810.340000 ;
        RECT 1705.940000 769.100000 1707.540000 810.340000 ;
        RECT 1622.940000 769.100000 1624.540000 810.340000 ;
        RECT 1622.940000 529.100000 1624.540000 630.040000 ;
        RECT 1814.780000 529.100000 1816.380000 630.040000 ;
        RECT 1705.940000 529.100000 1707.540000 630.040000 ;
        RECT 1705.940000 728.740000 1707.540000 772.300000 ;
        RECT 1814.780000 728.740000 1816.380000 772.300000 ;
        RECT 1897.780000 529.100000 1899.380000 630.040000 ;
        RECT 1897.780000 728.740000 1899.380000 772.300000 ;
        RECT 1814.780000 909.040000 1816.380000 952.300000 ;
        RECT 1705.940000 909.040000 1707.540000 952.300000 ;
        RECT 1622.940000 909.040000 1624.540000 952.300000 ;
        RECT 1897.780000 909.040000 1899.380000 952.300000 ;
        RECT 1039.100000 2038.300000 1042.300000 2055.100000 ;
        RECT 911.700000 1509.100000 913.300000 1580.780000 ;
        RECT 828.700000 1509.100000 830.300000 1580.780000 ;
        RECT 719.860000 1509.100000 721.460000 1580.780000 ;
        RECT 636.860000 1509.100000 638.460000 1580.780000 ;
        RECT 421.780000 1509.100000 423.380000 1580.780000 ;
        RECT 338.780000 1509.100000 340.380000 1580.780000 ;
        RECT 229.940000 1509.100000 231.540000 1580.780000 ;
        RECT 146.940000 1509.100000 148.540000 1580.780000 ;
        RECT 241.500000 1201.150000 243.100000 1262.300000 ;
        RECT 146.940000 1201.150000 148.540000 1262.300000 ;
        RECT 146.940000 1259.100000 148.540000 1282.750000 ;
        RECT 247.740000 1259.100000 249.340000 1282.750000 ;
        RECT 338.780000 1207.070000 340.380000 1262.300000 ;
        RECT 274.100000 1195.780000 279.300000 1197.380000 ;
        RECT 338.780000 1259.100000 340.380000 1282.750000 ;
        RECT 439.580000 1207.070000 441.180000 1262.300000 ;
        RECT 439.580000 1259.100000 441.180000 1282.750000 ;
        RECT 247.740000 1399.180000 249.340000 1432.300000 ;
        RECT 439.580000 1399.180000 441.180000 1432.300000 ;
        RECT 338.780000 1399.180000 340.380000 1432.300000 ;
        RECT 636.860000 1259.100000 638.460000 1282.750000 ;
        RECT 731.420000 1201.150000 733.020000 1262.300000 ;
        RECT 737.660000 1259.100000 739.260000 1282.750000 ;
        RECT 828.700000 1259.100000 830.300000 1282.750000 ;
        RECT 929.500000 1207.070000 931.100000 1262.300000 ;
        RECT 929.500000 1259.100000 931.100000 1282.750000 ;
        RECT 737.660000 1399.180000 739.260000 1432.300000 ;
        RECT 828.700000 1399.180000 830.300000 1432.300000 ;
        RECT 929.500000 1399.180000 931.100000 1432.300000 ;
        RECT 229.940000 1679.480000 231.540000 1752.300000 ;
        RECT 146.940000 1679.480000 148.540000 1752.300000 ;
        RECT 229.940000 1749.100000 231.540000 1761.080000 ;
        RECT 146.940000 1749.100000 148.540000 1761.080000 ;
        RECT 421.780000 1679.480000 423.380000 1752.300000 ;
        RECT 338.780000 1679.480000 340.380000 1752.300000 ;
        RECT 338.780000 1749.100000 340.380000 1761.080000 ;
        RECT 421.780000 1749.100000 423.380000 1761.080000 ;
        RECT 229.940000 1859.780000 231.540000 1912.300000 ;
        RECT 421.780000 1859.780000 423.380000 1912.300000 ;
        RECT 274.100000 2038.300000 277.300000 2055.100000 ;
        RECT 499.100000 2038.300000 502.300000 2055.100000 ;
        RECT 719.860000 1679.480000 721.460000 1752.300000 ;
        RECT 636.860000 1749.100000 638.460000 1761.080000 ;
        RECT 719.860000 1749.100000 721.460000 1761.080000 ;
        RECT 911.700000 1679.480000 913.300000 1752.300000 ;
        RECT 828.700000 1749.100000 830.300000 1761.080000 ;
        RECT 911.700000 1749.100000 913.300000 1761.080000 ;
        RECT 636.860000 1859.780000 638.460000 1912.300000 ;
        RECT 719.860000 1859.780000 721.460000 1912.300000 ;
        RECT 539.100000 2038.300000 542.300000 2055.100000 ;
        RECT 774.100000 2038.300000 777.300000 2055.100000 ;
        RECT 911.700000 1859.780000 913.300000 1912.300000 ;
        RECT 1009.100000 2038.300000 1012.300000 2055.100000 ;
        RECT 1407.860000 1509.100000 1409.460000 1592.620000 ;
        RECT 1324.860000 1509.100000 1326.460000 1592.620000 ;
        RECT 1209.780000 1509.100000 1211.380000 1592.620000 ;
        RECT 1126.780000 1509.100000 1128.380000 1592.620000 ;
        RECT 1897.780000 1509.100000 1899.380000 1580.780000 ;
        RECT 1814.780000 1509.100000 1816.380000 1580.780000 ;
        RECT 1705.940000 1509.100000 1707.540000 1580.780000 ;
        RECT 1622.940000 1509.100000 1624.540000 1580.780000 ;
        RECT 1126.780000 1259.100000 1128.380000 1294.590000 ;
        RECT 1227.580000 1212.990000 1229.180000 1262.300000 ;
        RECT 1227.580000 1259.100000 1229.180000 1294.590000 ;
        RECT 1425.660000 1212.990000 1427.260000 1262.300000 ;
        RECT 1324.860000 1259.100000 1326.460000 1294.590000 ;
        RECT 1425.660000 1259.100000 1427.260000 1294.590000 ;
        RECT 1227.580000 1411.020000 1229.180000 1432.300000 ;
        RECT 1324.860000 1411.020000 1326.460000 1432.300000 ;
        RECT 1425.660000 1411.020000 1427.260000 1432.300000 ;
        RECT 1622.940000 1259.100000 1624.540000 1282.750000 ;
        RECT 1717.500000 1201.150000 1719.100000 1262.300000 ;
        RECT 1723.740000 1259.100000 1725.340000 1282.750000 ;
        RECT 1814.780000 1259.100000 1816.380000 1282.750000 ;
        RECT 1915.580000 1207.070000 1917.180000 1262.300000 ;
        RECT 1915.580000 1259.100000 1917.180000 1282.750000 ;
        RECT 1723.740000 1399.180000 1725.340000 1432.300000 ;
        RECT 1622.940000 1399.180000 1624.540000 1432.300000 ;
        RECT 1915.580000 1399.180000 1917.180000 1432.300000 ;
        RECT 1126.780000 1749.100000 1128.380000 1772.920000 ;
        RECT 1126.780000 1691.320000 1128.380000 1752.300000 ;
        RECT 1209.780000 1749.100000 1211.380000 1772.920000 ;
        RECT 1209.780000 1691.320000 1211.380000 1752.300000 ;
        RECT 1407.860000 1749.100000 1409.460000 1772.920000 ;
        RECT 1324.860000 1749.100000 1326.460000 1772.920000 ;
        RECT 1324.860000 1691.320000 1326.460000 1752.300000 ;
        RECT 1407.860000 1691.320000 1409.460000 1752.300000 ;
        RECT 1209.780000 1871.620000 1211.380000 1912.300000 ;
        RECT 1274.100000 2038.300000 1277.300000 2055.100000 ;
        RECT 1324.860000 1871.620000 1326.460000 1912.300000 ;
        RECT 1407.860000 1871.620000 1409.460000 1912.300000 ;
        RECT 1519.100000 2038.300000 1522.300000 2055.100000 ;
        RECT 1539.100000 2038.300000 1542.300000 2055.100000 ;
        RECT 1705.940000 1679.480000 1707.540000 1752.300000 ;
        RECT 1622.940000 1749.100000 1624.540000 1761.080000 ;
        RECT 1705.940000 1749.100000 1707.540000 1761.080000 ;
        RECT 1814.780000 1749.100000 1816.380000 1761.080000 ;
        RECT 1897.780000 1679.480000 1899.380000 1752.300000 ;
        RECT 1897.780000 1749.100000 1899.380000 1761.080000 ;
        RECT 1622.940000 1859.780000 1624.540000 1912.300000 ;
        RECT 1814.780000 1859.780000 1816.380000 1912.300000 ;
        RECT 1705.940000 1859.780000 1707.540000 1912.300000 ;
        RECT 1774.100000 2038.300000 1777.300000 2055.100000 ;
        RECT 1897.780000 1859.780000 1899.380000 1912.300000 ;
        RECT 2029.100000 2038.300000 2032.300000 2055.100000 ;
        RECT 1039.100000 38.860000 1042.300000 39.340000 ;
        RECT 274.100000 38.860000 277.300000 39.340000 ;
        RECT 499.100000 38.860000 502.300000 39.340000 ;
        RECT 539.100000 38.860000 542.300000 39.340000 ;
        RECT 774.100000 38.860000 777.300000 39.340000 ;
        RECT 1009.100000 38.860000 1012.300000 39.340000 ;
        RECT 1274.100000 38.860000 1277.300000 39.340000 ;
        RECT 1519.100000 38.860000 1522.300000 39.340000 ;
        RECT 1539.100000 38.860000 1542.300000 39.340000 ;
        RECT 1774.100000 38.860000 1777.300000 39.340000 ;
        RECT 2029.100000 38.860000 2032.300000 39.340000 ;
        RECT 304.840000 245.040000 306.260000 246.640000 ;
        RECT 304.840000 1195.780000 306.260000 1197.380000 ;
      LAYER met5 ;
        RECT 0.000000 22.300000 2078.280000 33.500000 ;
        RECT 1039.100000 147.000000 1119.740000 148.600000 ;
        RECT 1039.100000 245.040000 1119.740000 246.640000 ;
        RECT 39.100000 279.100000 2039.180000 282.300000 ;
        RECT 1039.100000 345.030000 1119.740000 346.630000 ;
        RECT 1039.100000 443.070000 1119.740000 444.670000 ;
        RECT 39.100000 469.100000 2039.180000 472.300000 ;
        RECT 39.100000 529.100000 2039.180000 532.300000 ;
        RECT 1039.100000 643.180000 1119.740000 644.780000 ;
        RECT 1039.100000 724.140000 1119.740000 725.740000 ;
        RECT 39.100000 769.100000 2039.180000 772.300000 ;
        RECT 1039.100000 823.480000 1119.740000 825.080000 ;
        RECT 1039.100000 904.440000 1119.740000 906.040000 ;
        RECT 39.100000 949.100000 2039.180000 952.300000 ;
        RECT 39.100000 1019.100000 2039.180000 1022.300000 ;
        RECT 250.140000 147.000000 277.300000 148.600000 ;
        RECT 250.140000 241.710000 277.300000 243.310000 ;
        RECT 22.300000 147.000000 139.900000 148.600000 ;
        RECT 22.300000 241.710000 139.900000 243.310000 ;
        RECT 274.100000 147.000000 331.740000 148.600000 ;
        RECT 305.150000 245.040000 331.740000 246.640000 ;
        RECT 448.220000 147.000000 502.300000 148.600000 ;
        RECT 448.220000 245.040000 502.300000 246.640000 ;
        RECT 256.380000 339.110000 277.300000 340.710000 ;
        RECT 256.380000 437.150000 277.300000 438.750000 ;
        RECT 22.300000 339.110000 139.900000 340.710000 ;
        RECT 22.300000 279.100000 39.100000 282.300000 ;
        RECT 22.300000 437.150000 139.900000 438.750000 ;
        RECT 22.300000 469.100000 39.100000 472.300000 ;
        RECT 274.100000 339.110000 331.740000 340.710000 ;
        RECT 448.220000 339.110000 502.300000 340.710000 ;
        RECT 274.100000 437.150000 331.740000 438.750000 ;
        RECT 448.220000 437.150000 502.300000 438.750000 ;
        RECT 774.100000 147.000000 821.660000 148.600000 ;
        RECT 774.100000 245.040000 821.660000 246.640000 ;
        RECT 539.100000 147.000000 629.820000 148.600000 ;
        RECT 539.100000 241.710000 629.820000 243.310000 ;
        RECT 740.060000 147.000000 777.300000 148.600000 ;
        RECT 740.060000 241.710000 777.300000 243.310000 ;
        RECT 938.140000 147.000000 1012.300000 148.600000 ;
        RECT 938.140000 245.040000 1012.300000 246.640000 ;
        RECT 774.100000 339.110000 821.660000 340.710000 ;
        RECT 774.100000 437.150000 821.660000 438.750000 ;
        RECT 539.100000 339.110000 629.820000 340.710000 ;
        RECT 746.300000 339.110000 777.300000 340.710000 ;
        RECT 539.100000 437.150000 629.820000 438.750000 ;
        RECT 746.300000 437.150000 777.300000 438.750000 ;
        RECT 938.140000 339.110000 1012.300000 340.710000 ;
        RECT 938.140000 437.150000 1012.300000 438.750000 ;
        RECT 238.580000 637.260000 277.300000 638.860000 ;
        RECT 238.580000 718.220000 277.300000 719.820000 ;
        RECT 22.300000 637.260000 139.900000 638.860000 ;
        RECT 22.300000 529.100000 39.100000 532.300000 ;
        RECT 22.300000 718.220000 139.900000 719.820000 ;
        RECT 22.300000 769.100000 39.100000 772.300000 ;
        RECT 274.100000 637.260000 331.740000 638.860000 ;
        RECT 430.420000 637.260000 502.300000 638.860000 ;
        RECT 274.100000 718.220000 331.740000 719.820000 ;
        RECT 430.420000 718.220000 502.300000 719.820000 ;
        RECT 238.580000 817.560000 277.300000 819.160000 ;
        RECT 238.580000 898.520000 277.300000 900.120000 ;
        RECT 22.300000 817.560000 139.900000 819.160000 ;
        RECT 22.300000 898.520000 139.900000 900.120000 ;
        RECT 22.300000 949.100000 39.100000 952.300000 ;
        RECT 22.300000 1019.100000 39.100000 1022.300000 ;
        RECT 274.100000 817.560000 331.740000 819.160000 ;
        RECT 274.100000 898.520000 331.740000 900.120000 ;
        RECT 430.420000 817.560000 502.300000 819.160000 ;
        RECT 430.420000 898.520000 502.300000 900.120000 ;
        RECT 774.100000 637.260000 821.660000 638.860000 ;
        RECT 774.100000 718.220000 821.660000 719.820000 ;
        RECT 539.100000 637.260000 629.820000 638.860000 ;
        RECT 728.500000 637.260000 777.300000 638.860000 ;
        RECT 539.100000 718.220000 629.820000 719.820000 ;
        RECT 728.500000 718.220000 777.300000 719.820000 ;
        RECT 920.340000 637.260000 1012.300000 638.860000 ;
        RECT 920.340000 718.220000 1012.300000 719.820000 ;
        RECT 774.100000 817.560000 821.660000 819.160000 ;
        RECT 774.100000 898.520000 821.660000 900.120000 ;
        RECT 539.100000 817.560000 629.820000 819.160000 ;
        RECT 539.100000 898.520000 629.820000 900.120000 ;
        RECT 728.500000 817.560000 777.300000 819.160000 ;
        RECT 728.500000 898.520000 777.300000 900.120000 ;
        RECT 920.340000 817.560000 1012.300000 819.160000 ;
        RECT 920.340000 898.520000 1012.300000 900.120000 ;
        RECT 1539.100000 147.000000 1615.900000 148.600000 ;
        RECT 1539.100000 241.710000 1615.900000 243.310000 ;
        RECT 1539.100000 339.110000 1615.900000 340.710000 ;
        RECT 1539.100000 437.150000 1615.900000 438.750000 ;
        RECT 1274.100000 147.000000 1317.820000 148.600000 ;
        RECT 1274.100000 245.040000 1317.820000 246.640000 ;
        RECT 1236.220000 147.000000 1277.300000 148.600000 ;
        RECT 1236.220000 245.040000 1277.300000 246.640000 ;
        RECT 1434.300000 147.000000 1522.300000 148.600000 ;
        RECT 1434.300000 245.040000 1522.300000 246.640000 ;
        RECT 1274.100000 345.030000 1317.820000 346.630000 ;
        RECT 1274.100000 443.070000 1317.820000 444.670000 ;
        RECT 1236.220000 345.030000 1277.300000 346.630000 ;
        RECT 1236.220000 443.070000 1277.300000 444.670000 ;
        RECT 1434.300000 345.030000 1522.300000 346.630000 ;
        RECT 1434.300000 443.070000 1522.300000 444.670000 ;
        RECT 1726.140000 147.000000 1777.300000 148.600000 ;
        RECT 1774.100000 147.000000 1807.740000 148.600000 ;
        RECT 1726.140000 241.710000 1777.300000 243.310000 ;
        RECT 1774.100000 245.040000 1807.740000 246.640000 ;
        RECT 1924.220000 147.000000 2032.300000 148.600000 ;
        RECT 1924.220000 245.040000 2032.300000 246.640000 ;
        RECT 1732.380000 339.110000 1777.300000 340.710000 ;
        RECT 1774.100000 339.110000 1807.740000 340.710000 ;
        RECT 1732.380000 437.150000 1777.300000 438.750000 ;
        RECT 1774.100000 437.150000 1807.740000 438.750000 ;
        RECT 1924.220000 339.110000 2032.300000 340.710000 ;
        RECT 2039.180000 279.100000 2055.980000 282.300000 ;
        RECT 1924.220000 437.150000 2032.300000 438.750000 ;
        RECT 2039.180000 469.100000 2055.980000 472.300000 ;
        RECT 1539.100000 637.260000 1615.900000 638.860000 ;
        RECT 1539.100000 718.220000 1615.900000 719.820000 ;
        RECT 1539.100000 817.560000 1615.900000 819.160000 ;
        RECT 1539.100000 898.520000 1615.900000 900.120000 ;
        RECT 1274.100000 643.180000 1317.820000 644.780000 ;
        RECT 1274.100000 724.140000 1317.820000 725.740000 ;
        RECT 1218.420000 643.180000 1277.300000 644.780000 ;
        RECT 1218.420000 724.140000 1277.300000 725.740000 ;
        RECT 1416.500000 643.180000 1522.300000 644.780000 ;
        RECT 1416.500000 724.140000 1522.300000 725.740000 ;
        RECT 1274.100000 823.480000 1317.820000 825.080000 ;
        RECT 1274.100000 904.440000 1317.820000 906.040000 ;
        RECT 1218.420000 823.480000 1277.300000 825.080000 ;
        RECT 1218.420000 904.440000 1277.300000 906.040000 ;
        RECT 1416.500000 904.440000 1522.300000 906.040000 ;
        RECT 1416.500000 823.480000 1522.300000 825.080000 ;
        RECT 1714.580000 637.260000 1777.300000 638.860000 ;
        RECT 1774.100000 637.260000 1807.740000 638.860000 ;
        RECT 1714.580000 718.220000 1777.300000 719.820000 ;
        RECT 1774.100000 718.220000 1807.740000 719.820000 ;
        RECT 1906.420000 637.260000 2032.300000 638.860000 ;
        RECT 2039.180000 529.100000 2055.980000 532.300000 ;
        RECT 1906.420000 718.220000 2032.300000 719.820000 ;
        RECT 2039.180000 769.100000 2055.980000 772.300000 ;
        RECT 1714.580000 817.560000 1777.300000 819.160000 ;
        RECT 1774.100000 817.560000 1807.740000 819.160000 ;
        RECT 1714.580000 898.520000 1777.300000 900.120000 ;
        RECT 1774.100000 898.520000 1807.740000 900.120000 ;
        RECT 1906.420000 817.560000 2032.300000 819.160000 ;
        RECT 1906.420000 898.520000 2032.300000 900.120000 ;
        RECT 2039.180000 949.100000 2055.980000 952.300000 ;
        RECT 2039.180000 1019.100000 2055.980000 1022.300000 ;
        RECT 1039.100000 1103.660000 1119.740000 1105.260000 ;
        RECT 1039.100000 1201.700000 1119.740000 1203.300000 ;
        RECT 39.100000 1259.100000 2039.180000 1262.300000 ;
        RECT 1039.100000 1301.690000 1119.740000 1303.290000 ;
        RECT 1039.100000 1399.730000 1119.740000 1401.330000 ;
        RECT 39.100000 1429.100000 2039.180000 1432.300000 ;
        RECT 39.100000 1509.100000 2039.180000 1512.300000 ;
        RECT 1039.100000 1599.840000 1119.740000 1601.440000 ;
        RECT 1039.100000 1680.800000 1119.740000 1682.400000 ;
        RECT 39.100000 1749.100000 2039.180000 1752.300000 ;
        RECT 1039.100000 1780.140000 1119.740000 1781.740000 ;
        RECT 1039.100000 1861.100000 1119.740000 1862.700000 ;
        RECT 39.100000 1909.100000 2039.180000 1912.300000 ;
        RECT 39.100000 1999.100000 2039.180000 2002.300000 ;
        RECT 0.000000 2043.900000 2078.280000 2055.100000 ;
        RECT 250.140000 1097.740000 277.300000 1099.340000 ;
        RECT 256.380000 1289.850000 277.300000 1291.450000 ;
        RECT 250.140000 1192.450000 277.300000 1194.050000 ;
        RECT 22.300000 1097.740000 139.900000 1099.340000 ;
        RECT 22.300000 1289.850000 139.900000 1291.450000 ;
        RECT 22.300000 1192.450000 139.900000 1194.050000 ;
        RECT 22.300000 1259.100000 39.100000 1262.300000 ;
        RECT 274.100000 1097.740000 331.740000 1099.340000 ;
        RECT 448.220000 1097.740000 502.300000 1099.340000 ;
        RECT 305.150000 1195.780000 331.740000 1197.380000 ;
        RECT 274.100000 1289.850000 331.740000 1291.450000 ;
        RECT 448.220000 1195.780000 502.300000 1197.380000 ;
        RECT 448.220000 1289.850000 502.300000 1291.450000 ;
        RECT 256.380000 1387.890000 277.300000 1389.490000 ;
        RECT 22.300000 1387.890000 139.900000 1389.490000 ;
        RECT 22.300000 1429.100000 39.100000 1432.300000 ;
        RECT 22.300000 1509.100000 39.100000 1512.300000 ;
        RECT 274.100000 1387.890000 331.740000 1389.490000 ;
        RECT 448.220000 1387.890000 502.300000 1389.490000 ;
        RECT 774.100000 1097.740000 821.660000 1099.340000 ;
        RECT 774.100000 1195.780000 821.660000 1197.380000 ;
        RECT 774.100000 1289.850000 821.660000 1291.450000 ;
        RECT 539.100000 1097.740000 629.820000 1099.340000 ;
        RECT 740.060000 1097.740000 777.300000 1099.340000 ;
        RECT 539.100000 1192.450000 629.820000 1194.050000 ;
        RECT 539.100000 1289.850000 629.820000 1291.450000 ;
        RECT 740.060000 1192.450000 777.300000 1194.050000 ;
        RECT 746.300000 1289.850000 777.300000 1291.450000 ;
        RECT 938.140000 1097.740000 1012.300000 1099.340000 ;
        RECT 938.140000 1195.780000 1012.300000 1197.380000 ;
        RECT 938.140000 1289.850000 1012.300000 1291.450000 ;
        RECT 774.100000 1387.890000 821.660000 1389.490000 ;
        RECT 539.100000 1387.890000 629.820000 1389.490000 ;
        RECT 746.300000 1387.890000 777.300000 1389.490000 ;
        RECT 938.140000 1387.890000 1012.300000 1389.490000 ;
        RECT 238.580000 1588.000000 277.300000 1589.600000 ;
        RECT 238.580000 1668.960000 277.300000 1670.560000 ;
        RECT 238.580000 1768.300000 277.300000 1769.900000 ;
        RECT 22.300000 1588.000000 139.900000 1589.600000 ;
        RECT 22.300000 1668.960000 139.900000 1670.560000 ;
        RECT 22.300000 1768.300000 139.900000 1769.900000 ;
        RECT 22.300000 1749.100000 39.100000 1752.300000 ;
        RECT 274.100000 1588.000000 331.740000 1589.600000 ;
        RECT 274.100000 1668.960000 331.740000 1670.560000 ;
        RECT 430.420000 1588.000000 502.300000 1589.600000 ;
        RECT 430.420000 1668.960000 502.300000 1670.560000 ;
        RECT 274.100000 1768.300000 331.740000 1769.900000 ;
        RECT 430.420000 1768.300000 502.300000 1769.900000 ;
        RECT 238.580000 1849.260000 277.300000 1850.860000 ;
        RECT 22.300000 1849.260000 139.900000 1850.860000 ;
        RECT 22.300000 1909.100000 39.100000 1912.300000 ;
        RECT 22.300000 1999.100000 39.100000 2002.300000 ;
        RECT 274.100000 1849.260000 331.740000 1850.860000 ;
        RECT 430.420000 1849.260000 502.300000 1850.860000 ;
        RECT 774.100000 1588.000000 821.660000 1589.600000 ;
        RECT 774.100000 1668.960000 821.660000 1670.560000 ;
        RECT 774.100000 1768.300000 821.660000 1769.900000 ;
        RECT 539.100000 1588.000000 629.820000 1589.600000 ;
        RECT 539.100000 1668.960000 629.820000 1670.560000 ;
        RECT 728.500000 1588.000000 777.300000 1589.600000 ;
        RECT 728.500000 1668.960000 777.300000 1670.560000 ;
        RECT 539.100000 1768.300000 629.820000 1769.900000 ;
        RECT 728.500000 1768.300000 777.300000 1769.900000 ;
        RECT 920.340000 1588.000000 1012.300000 1589.600000 ;
        RECT 920.340000 1668.960000 1012.300000 1670.560000 ;
        RECT 920.340000 1768.300000 1012.300000 1769.900000 ;
        RECT 774.100000 1849.260000 821.660000 1850.860000 ;
        RECT 539.100000 1849.260000 629.820000 1850.860000 ;
        RECT 728.500000 1849.260000 777.300000 1850.860000 ;
        RECT 920.340000 1849.260000 1012.300000 1850.860000 ;
        RECT 1539.100000 1097.740000 1615.900000 1099.340000 ;
        RECT 1539.100000 1192.450000 1615.900000 1194.050000 ;
        RECT 1539.100000 1289.850000 1615.900000 1291.450000 ;
        RECT 1539.100000 1387.890000 1615.900000 1389.490000 ;
        RECT 1274.100000 1103.660000 1317.820000 1105.260000 ;
        RECT 1274.100000 1201.700000 1317.820000 1203.300000 ;
        RECT 1236.220000 1103.660000 1277.300000 1105.260000 ;
        RECT 1236.220000 1201.700000 1277.300000 1203.300000 ;
        RECT 1434.300000 1103.660000 1522.300000 1105.260000 ;
        RECT 1434.300000 1201.700000 1522.300000 1203.300000 ;
        RECT 1274.100000 1301.690000 1317.820000 1303.290000 ;
        RECT 1274.100000 1399.730000 1317.820000 1401.330000 ;
        RECT 1236.220000 1301.690000 1277.300000 1303.290000 ;
        RECT 1236.220000 1399.730000 1277.300000 1401.330000 ;
        RECT 1434.300000 1301.690000 1522.300000 1303.290000 ;
        RECT 1434.300000 1399.730000 1522.300000 1401.330000 ;
        RECT 1726.140000 1097.740000 1777.300000 1099.340000 ;
        RECT 1774.100000 1097.740000 1807.740000 1099.340000 ;
        RECT 1726.140000 1192.450000 1777.300000 1194.050000 ;
        RECT 1774.100000 1195.780000 1807.740000 1197.380000 ;
        RECT 1732.380000 1289.850000 1777.300000 1291.450000 ;
        RECT 1774.100000 1289.850000 1807.740000 1291.450000 ;
        RECT 1924.220000 1097.740000 2032.300000 1099.340000 ;
        RECT 1924.220000 1289.850000 2032.300000 1291.450000 ;
        RECT 1924.220000 1195.780000 2032.300000 1197.380000 ;
        RECT 2039.180000 1259.100000 2055.980000 1262.300000 ;
        RECT 1732.380000 1387.890000 1777.300000 1389.490000 ;
        RECT 1774.100000 1387.890000 1807.740000 1389.490000 ;
        RECT 1924.220000 1387.890000 2032.300000 1389.490000 ;
        RECT 2039.180000 1429.100000 2055.980000 1432.300000 ;
        RECT 2039.180000 1509.100000 2055.980000 1512.300000 ;
        RECT 1539.100000 1588.000000 1615.900000 1589.600000 ;
        RECT 1539.100000 1668.960000 1615.900000 1670.560000 ;
        RECT 1539.100000 1768.300000 1615.900000 1769.900000 ;
        RECT 1539.100000 1849.260000 1615.900000 1850.860000 ;
        RECT 1274.100000 1599.840000 1317.820000 1601.440000 ;
        RECT 1274.100000 1680.800000 1317.820000 1682.400000 ;
        RECT 1274.100000 1780.140000 1317.820000 1781.740000 ;
        RECT 1218.420000 1599.840000 1277.300000 1601.440000 ;
        RECT 1218.420000 1680.800000 1277.300000 1682.400000 ;
        RECT 1218.420000 1780.140000 1277.300000 1781.740000 ;
        RECT 1416.500000 1599.840000 1522.300000 1601.440000 ;
        RECT 1416.500000 1680.800000 1522.300000 1682.400000 ;
        RECT 1416.500000 1780.140000 1522.300000 1781.740000 ;
        RECT 1274.100000 1861.100000 1317.820000 1862.700000 ;
        RECT 1218.420000 1861.100000 1277.300000 1862.700000 ;
        RECT 1416.500000 1861.100000 1522.300000 1862.700000 ;
        RECT 1714.580000 1588.000000 1777.300000 1589.600000 ;
        RECT 1774.100000 1588.000000 1807.740000 1589.600000 ;
        RECT 1714.580000 1668.960000 1777.300000 1670.560000 ;
        RECT 1774.100000 1668.960000 1807.740000 1670.560000 ;
        RECT 1714.580000 1768.300000 1777.300000 1769.900000 ;
        RECT 1774.100000 1768.300000 1807.740000 1769.900000 ;
        RECT 1906.420000 1588.000000 2032.300000 1589.600000 ;
        RECT 1906.420000 1668.960000 2032.300000 1670.560000 ;
        RECT 1906.420000 1768.300000 2032.300000 1769.900000 ;
        RECT 2039.180000 1749.100000 2055.980000 1752.300000 ;
        RECT 1714.580000 1849.260000 1777.300000 1850.860000 ;
        RECT 1774.100000 1849.260000 1807.740000 1850.860000 ;
        RECT 1906.420000 1849.260000 2032.300000 1850.860000 ;
        RECT 2039.180000 1909.100000 2055.980000 1912.300000 ;
        RECT 2039.180000 1999.100000 2055.980000 2002.300000 ;
        RECT 304.840000 245.040000 306.260000 246.640000 ;
        RECT 304.840000 1195.780000 306.260000 1197.380000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2061.580000 2066.880000 2072.780000 2078.080000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.580000 0.000000 2072.780000 11.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.500000 2066.880000 16.700000 2078.080000 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.500000 0.000000 16.700000 11.200000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2067.080000 2060.700000 2078.280000 2071.900000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 2060.700000 11.200000 2071.900000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2067.080000 5.500000 2078.280000 16.700000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000000 5.500000 11.200000 16.700000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met4 ;
        RECT 1019.100000 39.100000 1022.300000 2038.300000 ;
        RECT 789.100000 39.100000 792.300000 2038.300000 ;
        RECT 544.100000 39.100000 547.300000 2038.300000 ;
        RECT 529.100000 39.100000 532.300000 2038.300000 ;
        RECT 299.100000 39.100000 302.300000 2038.300000 ;
        RECT 5.500000 0.000000 16.700000 2078.080000 ;
        RECT 1999.100000 39.100000 2002.300000 2038.300000 ;
        RECT 1769.100000 39.100000 1772.300000 2038.300000 ;
        RECT 1554.100000 39.100000 1557.300000 2038.300000 ;
        RECT 1509.100000 39.100000 1512.300000 2038.300000 ;
        RECT 1279.100000 39.100000 1282.300000 2038.300000 ;
        RECT 1049.100000 39.100000 1052.300000 2038.300000 ;
        RECT 2061.580000 0.000000 2072.780000 2078.080000 ;
        RECT 932.700000 448.440000 934.300000 522.300000 ;
        RECT 740.860000 448.440000 742.460000 522.300000 ;
        RECT 442.780000 448.440000 444.380000 522.300000 ;
        RECT 335.580000 448.440000 337.180000 522.300000 ;
        RECT 250.940000 448.440000 252.540000 522.300000 ;
        RECT 143.740000 448.440000 145.340000 522.300000 ;
        RECT 244.700000 250.410000 246.300000 272.300000 ;
        RECT 442.780000 256.330000 444.380000 272.300000 ;
        RECT 335.580000 256.330000 337.180000 272.300000 ;
        RECT 244.700000 5.500000 246.300000 139.900000 ;
        RECT 143.740000 5.500000 145.340000 139.900000 ;
        RECT 442.780000 5.500000 444.380000 139.900000 ;
        RECT 335.580000 5.500000 337.180000 139.900000 ;
        RECT 299.100000 5.500000 302.300000 39.100000 ;
        RECT 250.940000 269.100000 252.540000 332.010000 ;
        RECT 143.740000 269.100000 145.340000 332.010000 ;
        RECT 335.580000 269.100000 337.180000 332.010000 ;
        RECT 442.780000 269.100000 444.380000 332.010000 ;
        RECT 734.620000 250.410000 736.220000 272.300000 ;
        RECT 932.700000 256.330000 934.300000 272.300000 ;
        RECT 825.500000 256.330000 827.100000 272.300000 ;
        RECT 734.620000 5.500000 736.220000 139.900000 ;
        RECT 633.660000 5.500000 635.260000 139.900000 ;
        RECT 544.100000 5.500000 547.300000 39.100000 ;
        RECT 529.100000 5.500000 532.300000 39.100000 ;
        RECT 742.570000 244.910000 745.070000 246.510000 ;
        RECT 743.020000 245.710000 744.620000 247.890000 ;
        RECT 932.700000 5.500000 934.300000 139.900000 ;
        RECT 825.500000 5.500000 827.100000 139.900000 ;
        RECT 789.100000 5.500000 792.300000 39.100000 ;
        RECT 1019.100000 5.500000 1022.300000 39.100000 ;
        RECT 633.660000 269.100000 635.260000 332.010000 ;
        RECT 740.860000 269.100000 742.460000 332.010000 ;
        RECT 825.500000 269.100000 827.100000 332.010000 ;
        RECT 932.700000 269.100000 934.300000 332.010000 ;
        RECT 424.980000 749.100000 426.580000 810.340000 ;
        RECT 335.580000 749.100000 337.180000 810.340000 ;
        RECT 233.140000 749.100000 234.740000 810.340000 ;
        RECT 143.740000 749.100000 145.340000 810.340000 ;
        RECT 233.140000 539.100000 234.740000 630.040000 ;
        RECT 143.740000 539.100000 145.340000 630.040000 ;
        RECT 143.740000 728.740000 145.340000 752.300000 ;
        RECT 233.140000 728.740000 234.740000 752.300000 ;
        RECT 335.580000 539.100000 337.180000 630.040000 ;
        RECT 424.980000 539.100000 426.580000 630.040000 ;
        RECT 335.580000 728.740000 337.180000 752.300000 ;
        RECT 424.980000 728.740000 426.580000 752.300000 ;
        RECT 233.140000 909.040000 234.740000 1002.300000 ;
        RECT 143.740000 909.040000 145.340000 1002.300000 ;
        RECT 424.980000 909.040000 426.580000 1002.300000 ;
        RECT 335.580000 909.040000 337.180000 1002.300000 ;
        RECT 914.900000 749.100000 916.500000 810.340000 ;
        RECT 825.500000 749.100000 827.100000 810.340000 ;
        RECT 723.060000 749.100000 724.660000 810.340000 ;
        RECT 633.660000 749.100000 635.260000 810.340000 ;
        RECT 633.660000 539.100000 635.260000 630.040000 ;
        RECT 723.060000 539.100000 724.660000 630.040000 ;
        RECT 633.660000 728.740000 635.260000 752.300000 ;
        RECT 723.060000 728.740000 724.660000 752.300000 ;
        RECT 825.500000 539.100000 827.100000 630.040000 ;
        RECT 914.900000 539.100000 916.500000 630.040000 ;
        RECT 825.500000 728.740000 827.100000 752.300000 ;
        RECT 914.900000 728.740000 916.500000 752.300000 ;
        RECT 723.060000 909.040000 724.660000 1002.300000 ;
        RECT 914.900000 909.040000 916.500000 1002.300000 ;
        RECT 1918.780000 448.440000 1920.380000 522.300000 ;
        RECT 1726.940000 448.440000 1728.540000 522.300000 ;
        RECT 1619.740000 448.440000 1621.340000 522.300000 ;
        RECT 1428.860000 454.360000 1430.460000 522.300000 ;
        RECT 1230.780000 454.360000 1232.380000 522.300000 ;
        RECT 1428.860000 256.330000 1430.460000 272.300000 ;
        RECT 1321.660000 256.330000 1323.260000 272.300000 ;
        RECT 1230.780000 256.330000 1232.380000 272.300000 ;
        RECT 1230.780000 5.500000 1232.380000 139.900000 ;
        RECT 1123.580000 5.500000 1125.180000 139.900000 ;
        RECT 1049.100000 5.500000 1052.300000 39.100000 ;
        RECT 1279.100000 5.500000 1282.300000 39.100000 ;
        RECT 1428.860000 5.500000 1430.460000 139.900000 ;
        RECT 1321.660000 5.500000 1323.260000 139.900000 ;
        RECT 1554.100000 5.500000 1557.300000 39.100000 ;
        RECT 1509.100000 5.500000 1512.300000 39.100000 ;
        RECT 1123.580000 269.100000 1125.180000 337.930000 ;
        RECT 1230.780000 269.100000 1232.380000 337.930000 ;
        RECT 1321.660000 269.100000 1323.260000 337.930000 ;
        RECT 1428.860000 269.100000 1430.460000 337.930000 ;
        RECT 1720.700000 250.410000 1722.300000 272.300000 ;
        RECT 1619.740000 250.410000 1621.340000 272.300000 ;
        RECT 1918.780000 256.330000 1920.380000 272.300000 ;
        RECT 1811.580000 256.330000 1813.180000 272.300000 ;
        RECT 1811.580000 5.500000 1813.180000 139.900000 ;
        RECT 1720.700000 5.500000 1722.300000 139.900000 ;
        RECT 1619.740000 5.500000 1621.340000 139.900000 ;
        RECT 1769.100000 5.500000 1772.300000 39.100000 ;
        RECT 1918.780000 5.500000 1920.380000 139.900000 ;
        RECT 1999.100000 5.500000 2002.300000 39.100000 ;
        RECT 1619.740000 269.100000 1621.340000 332.010000 ;
        RECT 1811.580000 269.100000 1813.180000 332.010000 ;
        RECT 1726.940000 269.100000 1728.540000 332.010000 ;
        RECT 1918.780000 269.100000 1920.380000 332.010000 ;
        RECT 1411.060000 749.100000 1412.660000 816.260000 ;
        RECT 1321.660000 749.100000 1323.260000 816.260000 ;
        RECT 1212.980000 749.100000 1214.580000 816.260000 ;
        RECT 1123.580000 749.100000 1125.180000 816.260000 ;
        RECT 1123.580000 539.100000 1125.180000 635.960000 ;
        RECT 1212.980000 539.100000 1214.580000 635.960000 ;
        RECT 1123.580000 734.660000 1125.180000 752.300000 ;
        RECT 1212.980000 734.660000 1214.580000 752.300000 ;
        RECT 1411.060000 539.100000 1412.660000 635.960000 ;
        RECT 1321.660000 539.100000 1323.260000 635.960000 ;
        RECT 1321.660000 734.660000 1323.260000 752.300000 ;
        RECT 1411.060000 734.660000 1412.660000 752.300000 ;
        RECT 1212.980000 914.960000 1214.580000 1002.300000 ;
        RECT 1411.060000 914.960000 1412.660000 1002.300000 ;
        RECT 1321.660000 914.960000 1323.260000 1002.300000 ;
        RECT 1900.980000 749.100000 1902.580000 810.340000 ;
        RECT 1811.580000 749.100000 1813.180000 810.340000 ;
        RECT 1709.140000 749.100000 1710.740000 810.340000 ;
        RECT 1619.740000 749.100000 1621.340000 810.340000 ;
        RECT 1619.740000 539.100000 1621.340000 630.040000 ;
        RECT 1811.580000 539.100000 1813.180000 630.040000 ;
        RECT 1709.140000 539.100000 1710.740000 630.040000 ;
        RECT 1709.140000 728.740000 1710.740000 752.300000 ;
        RECT 1811.580000 728.740000 1813.180000 752.300000 ;
        RECT 1900.980000 539.100000 1902.580000 630.040000 ;
        RECT 1900.980000 728.740000 1902.580000 752.300000 ;
        RECT 1811.580000 909.040000 1813.180000 1002.300000 ;
        RECT 1709.140000 909.040000 1710.740000 1002.300000 ;
        RECT 1619.740000 909.040000 1621.340000 1002.300000 ;
        RECT 1900.980000 909.040000 1902.580000 1002.300000 ;
        RECT 914.900000 1539.100000 916.500000 1580.780000 ;
        RECT 825.500000 1539.100000 827.100000 1580.780000 ;
        RECT 723.060000 1539.100000 724.660000 1580.780000 ;
        RECT 633.660000 1539.100000 635.260000 1580.780000 ;
        RECT 424.980000 1539.100000 426.580000 1580.780000 ;
        RECT 335.580000 1539.100000 337.180000 1580.780000 ;
        RECT 233.140000 1539.100000 234.740000 1580.780000 ;
        RECT 143.740000 1539.100000 145.340000 1580.780000 ;
        RECT 143.740000 1039.100000 145.340000 1090.640000 ;
        RECT 244.700000 1039.100000 246.300000 1090.640000 ;
        RECT 250.940000 1229.100000 252.540000 1282.750000 ;
        RECT 143.740000 1229.100000 145.340000 1282.750000 ;
        RECT 143.740000 1201.150000 145.340000 1232.300000 ;
        RECT 244.700000 1201.150000 246.300000 1232.300000 ;
        RECT 335.580000 1039.100000 337.180000 1090.640000 ;
        RECT 442.780000 1039.100000 444.380000 1090.640000 ;
        RECT 335.580000 1229.100000 337.180000 1282.750000 ;
        RECT 335.580000 1207.070000 337.180000 1232.300000 ;
        RECT 442.780000 1229.100000 444.380000 1282.750000 ;
        RECT 442.780000 1207.070000 444.380000 1232.300000 ;
        RECT 250.940000 1399.180000 252.540000 1482.300000 ;
        RECT 143.740000 1399.180000 145.340000 1482.300000 ;
        RECT 442.780000 1399.180000 444.380000 1482.300000 ;
        RECT 633.660000 1039.100000 635.260000 1090.640000 ;
        RECT 734.620000 1039.100000 736.220000 1090.640000 ;
        RECT 633.660000 1229.100000 635.260000 1282.750000 ;
        RECT 740.860000 1229.100000 742.460000 1282.750000 ;
        RECT 734.620000 1201.150000 736.220000 1232.300000 ;
        RECT 825.500000 1039.100000 827.100000 1090.640000 ;
        RECT 932.700000 1039.100000 934.300000 1090.640000 ;
        RECT 825.500000 1229.100000 827.100000 1282.750000 ;
        RECT 825.500000 1207.070000 827.100000 1232.300000 ;
        RECT 932.700000 1229.100000 934.300000 1282.750000 ;
        RECT 932.700000 1207.070000 934.300000 1232.300000 ;
        RECT 740.860000 1399.180000 742.460000 1482.300000 ;
        RECT 932.700000 1399.180000 934.300000 1482.300000 ;
        RECT 825.500000 1399.180000 827.100000 1482.300000 ;
        RECT 233.140000 1679.480000 234.740000 1712.300000 ;
        RECT 143.740000 1679.480000 145.340000 1712.300000 ;
        RECT 233.140000 1709.100000 234.740000 1761.080000 ;
        RECT 143.740000 1709.100000 145.340000 1761.080000 ;
        RECT 424.980000 1679.480000 426.580000 1712.300000 ;
        RECT 335.580000 1679.480000 337.180000 1712.300000 ;
        RECT 335.580000 1709.100000 337.180000 1761.080000 ;
        RECT 424.980000 1709.100000 426.580000 1761.080000 ;
        RECT 233.140000 1859.780000 234.740000 1962.300000 ;
        RECT 143.740000 1859.780000 145.340000 1962.300000 ;
        RECT 424.980000 1859.780000 426.580000 1962.300000 ;
        RECT 335.580000 1859.780000 337.180000 1962.300000 ;
        RECT 299.100000 2038.300000 302.300000 2071.900000 ;
        RECT 723.060000 1679.480000 724.660000 1712.300000 ;
        RECT 633.660000 1709.100000 635.260000 1761.080000 ;
        RECT 723.060000 1709.100000 724.660000 1761.080000 ;
        RECT 914.900000 1679.480000 916.500000 1712.300000 ;
        RECT 825.500000 1679.480000 827.100000 1712.300000 ;
        RECT 825.500000 1709.100000 827.100000 1761.080000 ;
        RECT 914.900000 1709.100000 916.500000 1761.080000 ;
        RECT 723.060000 1859.780000 724.660000 1962.300000 ;
        RECT 633.660000 1859.780000 635.260000 1962.300000 ;
        RECT 529.100000 2038.300000 532.300000 2071.900000 ;
        RECT 544.100000 2038.300000 547.300000 2071.900000 ;
        RECT 914.900000 1859.780000 916.500000 1962.300000 ;
        RECT 789.100000 2038.300000 792.300000 2071.900000 ;
        RECT 1019.100000 2038.300000 1022.300000 2071.900000 ;
        RECT 1411.060000 1539.100000 1412.660000 1592.620000 ;
        RECT 1321.660000 1539.100000 1323.260000 1592.620000 ;
        RECT 1212.980000 1539.100000 1214.580000 1592.620000 ;
        RECT 1123.580000 1539.100000 1125.180000 1592.620000 ;
        RECT 1900.980000 1539.100000 1902.580000 1580.780000 ;
        RECT 1811.580000 1539.100000 1813.180000 1580.780000 ;
        RECT 1709.140000 1539.100000 1710.740000 1580.780000 ;
        RECT 1619.740000 1539.100000 1621.340000 1580.780000 ;
        RECT 1123.580000 1039.100000 1125.180000 1096.560000 ;
        RECT 1230.780000 1039.100000 1232.380000 1096.560000 ;
        RECT 1123.580000 1229.100000 1125.180000 1294.590000 ;
        RECT 1230.780000 1229.100000 1232.380000 1294.590000 ;
        RECT 1230.780000 1212.990000 1232.380000 1232.300000 ;
        RECT 1321.660000 1039.100000 1323.260000 1096.560000 ;
        RECT 1428.860000 1039.100000 1430.460000 1096.560000 ;
        RECT 1321.660000 1229.100000 1323.260000 1294.590000 ;
        RECT 1321.660000 1212.990000 1323.260000 1232.300000 ;
        RECT 1428.860000 1229.100000 1430.460000 1294.590000 ;
        RECT 1428.860000 1212.990000 1430.460000 1232.300000 ;
        RECT 1230.780000 1411.020000 1232.380000 1482.300000 ;
        RECT 1428.860000 1411.020000 1430.460000 1482.300000 ;
        RECT 1619.740000 1039.100000 1621.340000 1090.640000 ;
        RECT 1720.700000 1039.100000 1722.300000 1090.640000 ;
        RECT 1811.580000 1039.100000 1813.180000 1090.640000 ;
        RECT 1619.740000 1229.100000 1621.340000 1282.750000 ;
        RECT 1811.580000 1229.100000 1813.180000 1282.750000 ;
        RECT 1726.940000 1229.100000 1728.540000 1282.750000 ;
        RECT 1720.700000 1201.150000 1722.300000 1232.300000 ;
        RECT 1811.580000 1207.070000 1813.180000 1232.300000 ;
        RECT 1918.780000 1039.100000 1920.380000 1090.640000 ;
        RECT 1918.780000 1229.100000 1920.380000 1282.750000 ;
        RECT 1918.780000 1207.070000 1920.380000 1232.300000 ;
        RECT 1726.940000 1399.180000 1728.540000 1482.300000 ;
        RECT 1918.780000 1399.180000 1920.380000 1482.300000 ;
        RECT 1123.580000 1709.100000 1125.180000 1772.920000 ;
        RECT 1123.580000 1691.320000 1125.180000 1712.300000 ;
        RECT 1212.980000 1709.100000 1214.580000 1772.920000 ;
        RECT 1212.980000 1691.320000 1214.580000 1712.300000 ;
        RECT 1411.060000 1709.100000 1412.660000 1772.920000 ;
        RECT 1321.660000 1709.100000 1323.260000 1772.920000 ;
        RECT 1321.660000 1691.320000 1323.260000 1712.300000 ;
        RECT 1411.060000 1691.320000 1412.660000 1712.300000 ;
        RECT 1212.980000 1871.620000 1214.580000 1962.300000 ;
        RECT 1049.100000 2038.300000 1052.300000 2071.900000 ;
        RECT 1279.100000 2038.300000 1282.300000 2071.900000 ;
        RECT 1411.060000 1871.620000 1412.660000 1962.300000 ;
        RECT 1554.100000 2038.300000 1557.300000 2071.900000 ;
        RECT 1509.100000 2038.300000 1512.300000 2071.900000 ;
        RECT 1811.580000 1679.480000 1813.180000 1712.300000 ;
        RECT 1709.140000 1679.480000 1710.740000 1712.300000 ;
        RECT 1619.740000 1679.480000 1621.340000 1712.300000 ;
        RECT 1619.740000 1709.100000 1621.340000 1761.080000 ;
        RECT 1811.580000 1709.100000 1813.180000 1761.080000 ;
        RECT 1709.140000 1709.100000 1710.740000 1761.080000 ;
        RECT 1900.980000 1679.480000 1902.580000 1712.300000 ;
        RECT 1900.980000 1709.100000 1902.580000 1761.080000 ;
        RECT 1709.140000 1859.780000 1710.740000 1962.300000 ;
        RECT 1769.100000 2038.300000 1772.300000 2071.900000 ;
        RECT 1900.980000 1859.780000 1902.580000 1962.300000 ;
        RECT 1999.100000 2038.300000 2002.300000 2071.900000 ;
        RECT 743.020000 247.090000 744.620000 248.690000 ;
        RECT 1619.740000 749.015000 1621.340000 749.345000 ;
        RECT 299.100000 2038.060000 302.300000 2038.540000 ;
        RECT 544.100000 2038.060000 547.300000 2038.540000 ;
        RECT 529.100000 2038.060000 532.300000 2038.540000 ;
        RECT 789.100000 2038.060000 792.300000 2038.540000 ;
        RECT 1019.100000 2038.060000 1022.300000 2038.540000 ;
        RECT 1049.100000 2038.060000 1052.300000 2038.540000 ;
        RECT 1279.100000 2038.060000 1282.300000 2038.540000 ;
        RECT 1509.100000 2038.060000 1512.300000 2038.540000 ;
        RECT 1554.100000 2038.060000 1557.300000 2038.540000 ;
        RECT 1769.100000 2038.060000 1772.300000 2038.540000 ;
        RECT 1999.100000 2038.060000 2002.300000 2038.540000 ;
        RECT 768.890000 1195.650000 770.310000 1197.250000 ;
      LAYER met5 ;
        RECT 39.100000 519.100000 2039.180000 522.300000 ;
        RECT 0.000000 5.500000 2078.280000 16.700000 ;
        RECT 39.100000 269.100000 2039.180000 272.300000 ;
        RECT 39.100000 539.100000 2039.180000 542.300000 ;
        RECT 39.100000 749.100000 2039.180000 752.300000 ;
        RECT 39.100000 999.100000 2039.180000 1002.300000 ;
        RECT 5.500000 519.100000 39.100000 522.300000 ;
        RECT 448.220000 143.800000 532.300000 145.400000 ;
        RECT 448.220000 248.240000 532.300000 249.840000 ;
        RECT 448.220000 335.910000 532.300000 337.510000 ;
        RECT 448.220000 440.350000 532.300000 441.950000 ;
        RECT 250.140000 143.800000 302.300000 145.400000 ;
        RECT 250.140000 244.910000 302.300000 246.510000 ;
        RECT 5.500000 143.800000 139.900000 145.400000 ;
        RECT 5.500000 244.910000 139.900000 246.510000 ;
        RECT 299.100000 143.800000 331.740000 145.400000 ;
        RECT 299.100000 248.240000 331.740000 249.840000 ;
        RECT 256.380000 335.910000 302.300000 337.510000 ;
        RECT 256.380000 440.350000 302.300000 441.950000 ;
        RECT 5.500000 335.910000 139.900000 337.510000 ;
        RECT 5.500000 269.100000 39.100000 272.300000 ;
        RECT 5.500000 440.350000 139.900000 441.950000 ;
        RECT 299.100000 335.910000 331.740000 337.510000 ;
        RECT 299.100000 440.350000 331.740000 441.950000 ;
        RECT 740.060000 143.800000 792.300000 145.400000 ;
        RECT 544.100000 143.800000 629.820000 145.400000 ;
        RECT 544.100000 244.910000 629.820000 246.510000 ;
        RECT 740.060000 244.910000 743.820000 246.510000 ;
        RECT 789.100000 143.800000 821.660000 145.400000 ;
        RECT 789.100000 248.240000 821.660000 249.840000 ;
        RECT 938.140000 143.800000 1022.300000 145.400000 ;
        RECT 938.140000 248.240000 1022.300000 249.840000 ;
        RECT 746.300000 335.910000 792.300000 337.510000 ;
        RECT 746.300000 440.350000 792.300000 441.950000 ;
        RECT 544.100000 335.910000 629.820000 337.510000 ;
        RECT 544.100000 440.350000 629.820000 441.950000 ;
        RECT 789.100000 335.910000 821.660000 337.510000 ;
        RECT 938.140000 335.910000 1022.300000 337.510000 ;
        RECT 789.100000 440.350000 821.660000 441.950000 ;
        RECT 938.140000 440.350000 1022.300000 441.950000 ;
        RECT 430.420000 634.060000 532.300000 635.660000 ;
        RECT 430.420000 721.420000 532.300000 723.020000 ;
        RECT 430.420000 814.360000 532.300000 815.960000 ;
        RECT 430.420000 901.720000 532.300000 903.320000 ;
        RECT 238.580000 634.060000 302.300000 635.660000 ;
        RECT 238.580000 721.420000 302.300000 723.020000 ;
        RECT 5.500000 634.060000 139.900000 635.660000 ;
        RECT 5.500000 539.100000 39.100000 542.300000 ;
        RECT 5.500000 721.420000 139.900000 723.020000 ;
        RECT 5.500000 749.100000 39.100000 752.300000 ;
        RECT 299.100000 634.060000 331.740000 635.660000 ;
        RECT 299.100000 721.420000 331.740000 723.020000 ;
        RECT 238.580000 814.360000 302.300000 815.960000 ;
        RECT 238.580000 901.720000 302.300000 903.320000 ;
        RECT 5.500000 814.360000 139.900000 815.960000 ;
        RECT 5.500000 901.720000 139.900000 903.320000 ;
        RECT 5.500000 999.100000 39.100000 1002.300000 ;
        RECT 299.100000 814.360000 331.740000 815.960000 ;
        RECT 299.100000 901.720000 331.740000 903.320000 ;
        RECT 728.500000 634.060000 792.300000 635.660000 ;
        RECT 728.500000 721.420000 792.300000 723.020000 ;
        RECT 544.100000 634.060000 629.820000 635.660000 ;
        RECT 544.100000 721.420000 629.820000 723.020000 ;
        RECT 789.100000 634.060000 821.660000 635.660000 ;
        RECT 920.340000 634.060000 1022.300000 635.660000 ;
        RECT 789.100000 721.420000 821.660000 723.020000 ;
        RECT 920.340000 721.420000 1022.300000 723.020000 ;
        RECT 728.500000 814.360000 792.300000 815.960000 ;
        RECT 728.500000 901.720000 792.300000 903.320000 ;
        RECT 544.100000 814.360000 629.820000 815.960000 ;
        RECT 544.100000 901.720000 629.820000 903.320000 ;
        RECT 789.100000 814.360000 821.660000 815.960000 ;
        RECT 789.100000 901.720000 821.660000 903.320000 ;
        RECT 920.340000 814.360000 1022.300000 815.960000 ;
        RECT 920.340000 901.720000 1022.300000 903.320000 ;
        RECT 2039.180000 519.100000 2072.780000 522.300000 ;
        RECT 1554.100000 143.800000 1615.900000 145.400000 ;
        RECT 1554.100000 244.910000 1615.900000 246.510000 ;
        RECT 1554.100000 335.910000 1615.900000 337.510000 ;
        RECT 1554.100000 440.350000 1615.900000 441.950000 ;
        RECT 1279.100000 143.800000 1317.820000 145.400000 ;
        RECT 1279.100000 248.240000 1317.820000 249.840000 ;
        RECT 1049.100000 143.800000 1119.740000 145.400000 ;
        RECT 1049.100000 248.240000 1119.740000 249.840000 ;
        RECT 1236.220000 143.800000 1282.300000 145.400000 ;
        RECT 1236.220000 248.240000 1282.300000 249.840000 ;
        RECT 1434.300000 143.800000 1512.300000 145.400000 ;
        RECT 1434.300000 248.240000 1512.300000 249.840000 ;
        RECT 1279.100000 341.830000 1317.820000 343.430000 ;
        RECT 1279.100000 446.270000 1317.820000 447.870000 ;
        RECT 1049.100000 341.830000 1119.740000 343.430000 ;
        RECT 1236.220000 341.830000 1282.300000 343.430000 ;
        RECT 1049.100000 446.270000 1119.740000 447.870000 ;
        RECT 1236.220000 446.270000 1282.300000 447.870000 ;
        RECT 1434.300000 341.830000 1512.300000 343.430000 ;
        RECT 1434.300000 446.270000 1512.300000 447.870000 ;
        RECT 1726.140000 143.800000 1772.300000 145.400000 ;
        RECT 1769.100000 143.800000 1807.740000 145.400000 ;
        RECT 1726.140000 244.910000 1772.300000 246.510000 ;
        RECT 1769.100000 248.240000 1807.740000 249.840000 ;
        RECT 1924.220000 143.800000 2002.300000 145.400000 ;
        RECT 1924.220000 248.240000 2002.300000 249.840000 ;
        RECT 1732.380000 335.910000 1772.300000 337.510000 ;
        RECT 1769.100000 335.910000 1807.740000 337.510000 ;
        RECT 1732.380000 440.350000 1772.300000 441.950000 ;
        RECT 1769.100000 440.350000 1807.740000 441.950000 ;
        RECT 1924.220000 335.910000 2002.300000 337.510000 ;
        RECT 2039.180000 269.100000 2072.780000 272.300000 ;
        RECT 1924.220000 440.350000 2002.300000 441.950000 ;
        RECT 1554.100000 634.060000 1615.900000 635.660000 ;
        RECT 1554.100000 721.420000 1615.900000 723.020000 ;
        RECT 1554.100000 814.360000 1615.900000 815.960000 ;
        RECT 1554.100000 901.720000 1615.900000 903.320000 ;
        RECT 1279.100000 639.980000 1317.820000 641.580000 ;
        RECT 1279.100000 727.340000 1317.820000 728.940000 ;
        RECT 1049.100000 639.980000 1119.740000 641.580000 ;
        RECT 1218.420000 639.980000 1282.300000 641.580000 ;
        RECT 1049.100000 727.340000 1119.740000 728.940000 ;
        RECT 1218.420000 727.340000 1282.300000 728.940000 ;
        RECT 1416.500000 639.980000 1512.300000 641.580000 ;
        RECT 1416.500000 727.340000 1512.300000 728.940000 ;
        RECT 1279.100000 907.640000 1317.820000 909.240000 ;
        RECT 1279.100000 820.280000 1317.820000 821.880000 ;
        RECT 1049.100000 907.640000 1119.740000 909.240000 ;
        RECT 1218.420000 907.640000 1282.300000 909.240000 ;
        RECT 1049.100000 820.280000 1119.740000 821.880000 ;
        RECT 1218.420000 820.280000 1282.300000 821.880000 ;
        RECT 1416.500000 907.640000 1512.300000 909.240000 ;
        RECT 1416.500000 820.280000 1512.300000 821.880000 ;
        RECT 1714.580000 634.060000 1772.300000 635.660000 ;
        RECT 1769.100000 634.060000 1807.740000 635.660000 ;
        RECT 1714.580000 721.420000 1772.300000 723.020000 ;
        RECT 1769.100000 721.420000 1807.740000 723.020000 ;
        RECT 1906.420000 634.060000 2002.300000 635.660000 ;
        RECT 2039.180000 539.100000 2072.780000 542.300000 ;
        RECT 1906.420000 721.420000 2002.300000 723.020000 ;
        RECT 2039.180000 749.100000 2072.780000 752.300000 ;
        RECT 1714.580000 814.360000 1772.300000 815.960000 ;
        RECT 1769.100000 814.360000 1807.740000 815.960000 ;
        RECT 1714.580000 901.720000 1772.300000 903.320000 ;
        RECT 1769.100000 901.720000 1807.740000 903.320000 ;
        RECT 1906.420000 814.360000 2002.300000 815.960000 ;
        RECT 1906.420000 901.720000 2002.300000 903.320000 ;
        RECT 2039.180000 999.100000 2072.780000 1002.300000 ;
        RECT 39.100000 1039.100000 2039.180000 1042.300000 ;
        RECT 39.100000 1229.100000 2039.180000 1232.300000 ;
        RECT 39.100000 1479.100000 2039.180000 1482.300000 ;
        RECT 39.100000 1539.100000 2039.180000 1542.300000 ;
        RECT 39.100000 1709.100000 2039.180000 1712.300000 ;
        RECT 39.100000 1959.100000 2039.180000 1962.300000 ;
        RECT 0.000000 2060.700000 2078.280000 2071.900000 ;
        RECT 448.220000 1094.540000 532.300000 1096.140000 ;
        RECT 448.220000 1286.650000 532.300000 1288.250000 ;
        RECT 448.220000 1198.980000 532.300000 1200.580000 ;
        RECT 448.220000 1391.090000 532.300000 1392.690000 ;
        RECT 250.140000 1094.540000 302.300000 1096.140000 ;
        RECT 250.140000 1195.650000 302.300000 1197.250000 ;
        RECT 256.380000 1286.650000 302.300000 1288.250000 ;
        RECT 5.500000 1094.540000 139.900000 1096.140000 ;
        RECT 5.500000 1039.100000 39.100000 1042.300000 ;
        RECT 5.500000 1286.650000 139.900000 1288.250000 ;
        RECT 5.500000 1195.650000 139.900000 1197.250000 ;
        RECT 5.500000 1229.100000 39.100000 1232.300000 ;
        RECT 299.100000 1094.540000 331.740000 1096.140000 ;
        RECT 299.100000 1198.980000 331.740000 1200.580000 ;
        RECT 299.100000 1286.650000 331.740000 1288.250000 ;
        RECT 256.380000 1391.090000 302.300000 1392.690000 ;
        RECT 5.500000 1391.090000 139.900000 1392.690000 ;
        RECT 5.500000 1479.100000 39.100000 1482.300000 ;
        RECT 5.500000 1539.100000 39.100000 1542.300000 ;
        RECT 299.100000 1391.090000 331.740000 1392.690000 ;
        RECT 740.060000 1094.540000 792.300000 1096.140000 ;
        RECT 746.300000 1286.650000 792.300000 1288.250000 ;
        RECT 544.100000 1094.540000 629.820000 1096.140000 ;
        RECT 544.100000 1195.650000 629.820000 1197.250000 ;
        RECT 544.100000 1286.650000 629.820000 1288.250000 ;
        RECT 740.060000 1195.650000 770.000000 1197.250000 ;
        RECT 789.100000 1094.540000 821.660000 1096.140000 ;
        RECT 938.140000 1094.540000 1022.300000 1096.140000 ;
        RECT 789.100000 1198.980000 821.660000 1200.580000 ;
        RECT 789.100000 1286.650000 821.660000 1288.250000 ;
        RECT 938.140000 1198.980000 1022.300000 1200.580000 ;
        RECT 938.140000 1286.650000 1022.300000 1288.250000 ;
        RECT 746.300000 1391.090000 792.300000 1392.690000 ;
        RECT 544.100000 1391.090000 629.820000 1392.690000 ;
        RECT 789.100000 1391.090000 821.660000 1392.690000 ;
        RECT 938.140000 1391.090000 1022.300000 1392.690000 ;
        RECT 430.420000 1584.800000 532.300000 1586.400000 ;
        RECT 430.420000 1672.160000 532.300000 1673.760000 ;
        RECT 430.420000 1765.100000 532.300000 1766.700000 ;
        RECT 430.420000 1852.460000 532.300000 1854.060000 ;
        RECT 238.580000 1584.800000 302.300000 1586.400000 ;
        RECT 238.580000 1672.160000 302.300000 1673.760000 ;
        RECT 238.580000 1765.100000 302.300000 1766.700000 ;
        RECT 5.500000 1584.800000 139.900000 1586.400000 ;
        RECT 5.500000 1672.160000 139.900000 1673.760000 ;
        RECT 5.500000 1765.100000 139.900000 1766.700000 ;
        RECT 5.500000 1709.100000 39.100000 1712.300000 ;
        RECT 299.100000 1584.800000 331.740000 1586.400000 ;
        RECT 299.100000 1672.160000 331.740000 1673.760000 ;
        RECT 299.100000 1765.100000 331.740000 1766.700000 ;
        RECT 238.580000 1852.460000 302.300000 1854.060000 ;
        RECT 5.500000 1852.460000 139.900000 1854.060000 ;
        RECT 5.500000 1959.100000 39.100000 1962.300000 ;
        RECT 299.100000 1852.460000 331.740000 1854.060000 ;
        RECT 728.500000 1584.800000 792.300000 1586.400000 ;
        RECT 728.500000 1672.160000 792.300000 1673.760000 ;
        RECT 728.500000 1765.100000 792.300000 1766.700000 ;
        RECT 544.100000 1584.800000 629.820000 1586.400000 ;
        RECT 544.100000 1672.160000 629.820000 1673.760000 ;
        RECT 544.100000 1765.100000 629.820000 1766.700000 ;
        RECT 789.100000 1584.800000 821.660000 1586.400000 ;
        RECT 789.100000 1672.160000 821.660000 1673.760000 ;
        RECT 920.340000 1584.800000 1022.300000 1586.400000 ;
        RECT 920.340000 1672.160000 1022.300000 1673.760000 ;
        RECT 789.100000 1765.100000 821.660000 1766.700000 ;
        RECT 920.340000 1765.100000 1022.300000 1766.700000 ;
        RECT 728.500000 1852.460000 792.300000 1854.060000 ;
        RECT 544.100000 1852.460000 629.820000 1854.060000 ;
        RECT 789.100000 1852.460000 821.660000 1854.060000 ;
        RECT 920.340000 1852.460000 1022.300000 1854.060000 ;
        RECT 1554.100000 1094.540000 1615.900000 1096.140000 ;
        RECT 1554.100000 1286.650000 1615.900000 1288.250000 ;
        RECT 1554.100000 1195.650000 1615.900000 1197.250000 ;
        RECT 1554.100000 1391.090000 1615.900000 1392.690000 ;
        RECT 1434.300000 1298.490000 1512.300000 1300.090000 ;
        RECT 1049.100000 1298.490000 1119.740000 1300.090000 ;
        RECT 1236.220000 1298.490000 1282.300000 1300.090000 ;
        RECT 1279.100000 1298.490000 1317.820000 1300.090000 ;
        RECT 1279.100000 1100.460000 1317.820000 1102.060000 ;
        RECT 1279.100000 1204.900000 1317.820000 1206.500000 ;
        RECT 1049.100000 1100.460000 1119.740000 1102.060000 ;
        RECT 1236.220000 1100.460000 1282.300000 1102.060000 ;
        RECT 1049.100000 1204.900000 1119.740000 1206.500000 ;
        RECT 1236.220000 1204.900000 1282.300000 1206.500000 ;
        RECT 1434.300000 1100.460000 1512.300000 1102.060000 ;
        RECT 1434.300000 1204.900000 1512.300000 1206.500000 ;
        RECT 1279.100000 1402.930000 1317.820000 1404.530000 ;
        RECT 1049.100000 1402.930000 1119.740000 1404.530000 ;
        RECT 1236.220000 1402.930000 1282.300000 1404.530000 ;
        RECT 1434.300000 1402.930000 1512.300000 1404.530000 ;
        RECT 1726.140000 1094.540000 1772.300000 1096.140000 ;
        RECT 1769.100000 1094.540000 1807.740000 1096.140000 ;
        RECT 1726.140000 1195.650000 1772.300000 1197.250000 ;
        RECT 1769.100000 1198.980000 1807.740000 1200.580000 ;
        RECT 1732.380000 1286.650000 1772.300000 1288.250000 ;
        RECT 1769.100000 1286.650000 1807.740000 1288.250000 ;
        RECT 1924.220000 1094.540000 2002.300000 1096.140000 ;
        RECT 2039.180000 1039.100000 2072.780000 1042.300000 ;
        RECT 1924.220000 1286.650000 2002.300000 1288.250000 ;
        RECT 1924.220000 1198.980000 2002.300000 1200.580000 ;
        RECT 2039.180000 1229.100000 2072.780000 1232.300000 ;
        RECT 1732.380000 1391.090000 1772.300000 1392.690000 ;
        RECT 1769.100000 1391.090000 1807.740000 1392.690000 ;
        RECT 1924.220000 1391.090000 2002.300000 1392.690000 ;
        RECT 2039.180000 1479.100000 2072.780000 1482.300000 ;
        RECT 2039.180000 1539.100000 2072.780000 1542.300000 ;
        RECT 1554.100000 1584.800000 1615.900000 1586.400000 ;
        RECT 1554.100000 1672.160000 1615.900000 1673.760000 ;
        RECT 1554.100000 1765.100000 1615.900000 1766.700000 ;
        RECT 1554.100000 1852.460000 1615.900000 1854.060000 ;
        RECT 1279.100000 1596.640000 1317.820000 1598.240000 ;
        RECT 1279.100000 1684.000000 1317.820000 1685.600000 ;
        RECT 1279.100000 1776.940000 1317.820000 1778.540000 ;
        RECT 1049.100000 1596.640000 1119.740000 1598.240000 ;
        RECT 1049.100000 1684.000000 1119.740000 1685.600000 ;
        RECT 1218.420000 1596.640000 1282.300000 1598.240000 ;
        RECT 1218.420000 1684.000000 1282.300000 1685.600000 ;
        RECT 1049.100000 1776.940000 1119.740000 1778.540000 ;
        RECT 1218.420000 1776.940000 1282.300000 1778.540000 ;
        RECT 1416.500000 1684.000000 1512.300000 1685.600000 ;
        RECT 1416.500000 1596.640000 1512.300000 1598.240000 ;
        RECT 1416.500000 1776.940000 1512.300000 1778.540000 ;
        RECT 1279.100000 1864.300000 1317.820000 1865.900000 ;
        RECT 1049.100000 1864.300000 1119.740000 1865.900000 ;
        RECT 1218.420000 1864.300000 1282.300000 1865.900000 ;
        RECT 1416.500000 1864.300000 1512.300000 1865.900000 ;
        RECT 1714.580000 1584.800000 1772.300000 1586.400000 ;
        RECT 1769.100000 1584.800000 1807.740000 1586.400000 ;
        RECT 1714.580000 1672.160000 1772.300000 1673.760000 ;
        RECT 1769.100000 1672.160000 1807.740000 1673.760000 ;
        RECT 1714.580000 1765.100000 1772.300000 1766.700000 ;
        RECT 1769.100000 1765.100000 1807.740000 1766.700000 ;
        RECT 1906.420000 1584.800000 2002.300000 1586.400000 ;
        RECT 1906.420000 1672.160000 2002.300000 1673.760000 ;
        RECT 1906.420000 1765.100000 2002.300000 1766.700000 ;
        RECT 2039.180000 1709.100000 2072.780000 1712.300000 ;
        RECT 1714.580000 1852.460000 1772.300000 1854.060000 ;
        RECT 1769.100000 1852.460000 1807.740000 1854.060000 ;
        RECT 1906.420000 1852.460000 2002.300000 1854.060000 ;
        RECT 2039.180000 1959.100000 2072.780000 1962.300000 ;
        RECT 742.570000 244.910000 745.070000 246.510000 ;
        RECT 768.890000 1195.650000 770.310000 1197.250000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2078.280000 2078.080000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2078.280000 2078.080000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 2078.280000 2078.080000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 2078.280000 2078.080000 ;
    LAYER met4 ;
      RECT 0.000000 0.000000 2078.280000 2078.080000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2078.280000 2078.080000 ;
  END
END temp_wrapper

END LIBRARY
