##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Fri Dec 11 23:33:41 2020
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ldo
  CLASS BLOCK ;
  SIZE 311.040000 BY 311.540000 ;
  FOREIGN ldo 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.528 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.479 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 85.8669 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 461.144 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 98.28 LAYER met3  ;
    ANTENNAMAXAREACAR 8.7355 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.1293 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.171002 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 155.210000 0.000000 155.350000 0.485000 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.185 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.25 LAYER met2  ;
    ANTENNAMAXAREACAR 5.88529 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.1293 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.0834667 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 57.8805 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 313.376 LAYER met3  ;
    ANTENNAGATEAREA 50.88 LAYER met3  ;
    ANTENNAMAXAREACAR 18.0309 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 88.0698 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.312857 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 156.170000 0.000000 156.310000 0.485000 ;
    END
  END reset
  PIN mode_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.718 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.67 LAYER met2  ;
    ANTENNAMAXAREACAR 6.72633 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.5399 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.122381 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 187.850000 311.055000 187.990000 311.540000 ;
    END
  END mode_sel[1]
  PIN mode_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.8432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.42 LAYER met2  ;
    ANTENNAMAXAREACAR 29.4888 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 145.261 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.122381 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 180.170000 311.055000 180.310000 311.540000 ;
    END
  END mode_sel[0]
  PIN std_ctrl_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.491 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.125 LAYER met2  ;
    ANTENNAMAXAREACAR 8.23351 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.9871 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0456889 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 185.450000 311.055000 185.590000 311.540000 ;
    END
  END std_ctrl_in
  PIN std_pt_in_cnt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.8126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.729 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.09 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4272 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.9829 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.122381 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 136.010000 311.055000 136.150000 311.540000 ;
    END
  END std_pt_in_cnt[8]
  PIN std_pt_in_cnt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 109.2 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.67 LAYER met2  ;
    ANTENNAMAXAREACAR 9.32319 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.1093 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0833726 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 131.690000 311.055000 131.830000 311.540000 ;
    END
  END std_pt_in_cnt[7]
  PIN std_pt_in_cnt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.2214 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.537 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.92 LAYER met2  ;
    ANTENNAMAXAREACAR 6.48743 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.5531 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0979357 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 132.650000 311.055000 132.790000 311.540000 ;
    END
  END std_pt_in_cnt[6]
  PIN std_pt_in_cnt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0363 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.1735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.3834 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.875 LAYER met3  ;
    ANTENNAMAXAREACAR 8.18312 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 41.4577 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.143467 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 151.075000 0.595000 151.215000 ;
    END
  END std_pt_in_cnt[5]
  PIN std_pt_in_cnt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3915 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8495 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 41.4348 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 221.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.17 LAYER met3  ;
    ANTENNAMAXAREACAR 9.26564 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 46.1904 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.133539 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 0.000000 147.745000 0.595000 147.885000 ;
    END
  END std_pt_in_cnt[4]
  PIN std_pt_in_cnt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2127 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9555 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 62.8824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 338.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 12.375 LAYER met3  ;
    ANTENNAMAXAREACAR 8.81038 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.0597 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.207911 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 310.445000 138.495000 311.040000 138.635000 ;
    END
  END std_pt_in_cnt[3]
  PIN std_pt_in_cnt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1127 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.4555 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.38345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.125 LAYER met2  ;
    ANTENNAMAXAREACAR 3.01911 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.2627 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.1768 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.288 LAYER met3  ;
    ANTENNAGATEAREA 9 LAYER met3  ;
    ANTENNAMAXAREACAR 7.96252 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 39.3538 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.243467 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 310.445000 162.915000 311.040000 163.055000 ;
    END
  END std_pt_in_cnt[2]
  PIN std_pt_in_cnt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3471 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4983 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.3776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 216.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 6.75 LAYER met3  ;
    ANTENNAMAXAREACAR 8.94978 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 45.6131 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.1368 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 310.445000 157.365000 311.040000 157.505000 ;
    END
  END std_pt_in_cnt[1]
  PIN std_pt_in_cnt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4803 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.6315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.2365 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.375 LAYER met2  ;
    ANTENNAMAXAREACAR 3.30163 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.1881 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.0775407 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.3098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.456 LAYER met3  ;
    ANTENNAGATEAREA 4.5 LAYER met3  ;
    ANTENNAMAXAREACAR 3.5927 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 16.845 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0812444 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 310.445000 165.505000 311.040000 165.645000 ;
    END
  END std_pt_in_cnt[0]
  PIN cmp_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.1965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 36.5355 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 195.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.125 LAYER met3  ;
    ANTENNAMAXAREACAR 32.8116 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.213 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0812444 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 310.445000 139.235000 311.040000 139.375000 ;
    END
  END cmp_out
  PIN ctrl_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.59625 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.8826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 89.089 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.625 LAYER met2  ;
    ANTENNAMAXAREACAR 3.88337 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.4723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0456889 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 140.810000 311.055000 140.950000 311.540000 ;
    END
  END ctrl_out[8]
  PIN ctrl_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.59625 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.1548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.988 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.17 LAYER met2  ;
    ANTENNAMAXAREACAR 4.55587 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.7351 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.122381 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 130.730000 311.055000 130.870000 311.540000 ;
    END
  END ctrl_out[7]
  PIN ctrl_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.64125 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.9908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.728 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.125 LAYER met2  ;
    ANTENNAMAXAREACAR 15.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.2049 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0456889 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 120.650000 311.055000 120.790000 311.540000 ;
    END
  END ctrl_out[6]
  PIN ctrl_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.9607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.6425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.59625 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.0586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.44 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.17 LAYER met3  ;
    ANTENNAMAXAREACAR 3.73856 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 18.6177 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.0853666 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 119.690000 311.055000 119.830000 311.540000 ;
    END
  END ctrl_out[5]
  PIN ctrl_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.64125 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.6866 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 98.217 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.125 LAYER met2  ;
    ANTENNAMAXAREACAR 17.8816 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.8902 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0456889 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 152.330000 311.055000 152.470000 311.540000 ;
    END
  END ctrl_out[4]
  PIN ctrl_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.59625 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.17 LAYER met2  ;
    ANTENNAMAXAREACAR 3.85907 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.521 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0856635 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 163.370000 311.055000 163.510000 311.540000 ;
    END
  END ctrl_out[3]
  PIN ctrl_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.59625 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.0924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.17 LAYER met2  ;
    ANTENNAMAXAREACAR 3.62969 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0772365 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 173.450000 311.055000 173.590000 311.540000 ;
    END
  END ctrl_out[2]
  PIN ctrl_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.64125 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.978 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.5 LAYER met2  ;
    ANTENNAMAXAREACAR 5.13738 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.5091 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0456889 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 186.410000 311.055000 186.550000 311.540000 ;
    END
  END ctrl_out[1]
  PIN ctrl_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.59625 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.5012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.838 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 9.42 LAYER met2  ;
    ANTENNAMAXAREACAR 3.26455 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.1492 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.122381 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 188.810000 311.055000 188.950000 311.540000 ;
    END
  END ctrl_out[0]
  PIN VREF
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0804 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.3345 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 310.445000 76.705000 311.040000 76.845000 ;
    END
  END VREF
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.400000 309.740000 16.200000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.200000 309.740000 27.000000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.000000 309.740000 37.800000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.800000 309.740000 48.600000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.600000 309.740000 59.400000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.400000 309.740000 70.200000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.200000 309.740000 81.000000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.000000 309.740000 91.800000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.800000 309.740000 102.600000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.600000 309.740000 113.400000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.400000 309.740000 124.200000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 133.200000 309.740000 135.000000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.000000 309.740000 145.800000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.800000 309.740000 156.600000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.600000 309.740000 167.400000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 176.400000 309.740000 178.200000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 187.200000 309.740000 189.000000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 198.000000 309.740000 199.800000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.800000 309.740000 210.600000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.600000 309.740000 221.400000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 230.400000 309.740000 232.200000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 241.200000 309.740000 243.000000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 252.000000 309.740000 253.800000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 262.800000 309.740000 264.600000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 273.600000 309.740000 275.400000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.400000 309.740000 286.200000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 295.200000 309.740000 297.000000 311.540000 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.040000 304.100000 311.040000 306.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 304.100000 2.000000 306.100000 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.040000 4.330000 311.040000 6.330000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 4.330000 2.000000 6.330000 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.880000 309.540000 306.880000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.880000 0.000000 306.880000 2.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.160000 309.540000 6.160000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.160000 0.000000 6.160000 2.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 154.800000 75.225000 156.600000 76.475000 ;
        RECT 154.800000 115.925000 156.600000 117.175000 ;
        RECT 154.800000 83.365000 156.600000 84.615000 ;
        RECT 154.800000 91.505000 156.600000 92.755000 ;
        RECT 154.800000 99.645000 156.600000 100.895000 ;
        RECT 154.800000 107.785000 156.600000 109.035000 ;
        RECT 154.800000 124.065000 156.600000 125.315000 ;
        RECT 154.800000 132.205000 156.600000 133.455000 ;
        RECT 154.800000 140.345000 156.600000 141.595000 ;
        RECT 154.800000 148.485000 156.600000 149.735000 ;
        RECT 4.160000 18.245000 6.160000 19.495000 ;
        RECT 4.160000 10.615000 6.160000 11.355000 ;
        RECT 4.160000 34.525000 6.160000 35.775000 ;
        RECT 4.160000 26.385000 6.160000 27.635000 ;
        RECT 4.160000 50.805000 6.160000 52.055000 ;
        RECT 4.160000 42.665000 6.160000 43.915000 ;
        RECT 4.160000 75.225000 6.160000 76.475000 ;
        RECT 4.160000 67.085000 6.160000 68.335000 ;
        RECT 4.160000 58.945000 6.160000 60.195000 ;
        RECT 14.400000 75.225000 16.200000 76.475000 ;
        RECT 25.200000 75.225000 27.000000 76.475000 ;
        RECT 36.000000 75.225000 37.800000 76.475000 ;
        RECT 57.600000 75.225000 59.400000 76.475000 ;
        RECT 46.800000 75.225000 48.600000 76.475000 ;
        RECT 68.400000 75.225000 70.200000 76.475000 ;
        RECT 90.000000 75.225000 91.800000 76.475000 ;
        RECT 79.200000 75.225000 81.000000 76.475000 ;
        RECT 111.600000 75.225000 113.400000 76.475000 ;
        RECT 100.800000 75.225000 102.600000 76.475000 ;
        RECT 133.200000 75.225000 135.000000 76.475000 ;
        RECT 122.400000 75.225000 124.200000 76.475000 ;
        RECT 144.000000 75.225000 145.800000 76.475000 ;
        RECT 68.400000 115.925000 70.200000 117.175000 ;
        RECT 57.600000 115.925000 59.400000 117.175000 ;
        RECT 46.800000 115.925000 48.600000 117.175000 ;
        RECT 36.000000 115.925000 37.800000 117.175000 ;
        RECT 25.200000 115.925000 27.000000 117.175000 ;
        RECT 14.400000 115.925000 16.200000 117.175000 ;
        RECT 4.160000 115.925000 6.160000 117.175000 ;
        RECT 4.160000 83.365000 6.160000 84.615000 ;
        RECT 14.400000 83.365000 16.200000 84.615000 ;
        RECT 4.160000 91.505000 6.160000 92.755000 ;
        RECT 14.400000 91.505000 16.200000 92.755000 ;
        RECT 36.000000 83.365000 37.800000 84.615000 ;
        RECT 25.200000 83.365000 27.000000 84.615000 ;
        RECT 36.000000 91.505000 37.800000 92.755000 ;
        RECT 25.200000 91.505000 27.000000 92.755000 ;
        RECT 14.400000 107.785000 16.200000 109.035000 ;
        RECT 14.400000 99.645000 16.200000 100.895000 ;
        RECT 4.160000 107.785000 6.160000 109.035000 ;
        RECT 4.160000 99.645000 6.160000 100.895000 ;
        RECT 25.200000 99.645000 27.000000 100.895000 ;
        RECT 25.200000 107.785000 27.000000 109.035000 ;
        RECT 36.000000 99.645000 37.800000 100.895000 ;
        RECT 36.000000 107.785000 37.800000 109.035000 ;
        RECT 57.600000 83.365000 59.400000 84.615000 ;
        RECT 57.600000 91.505000 59.400000 92.755000 ;
        RECT 46.800000 91.505000 48.600000 92.755000 ;
        RECT 46.800000 83.365000 48.600000 84.615000 ;
        RECT 68.400000 91.505000 70.200000 92.755000 ;
        RECT 68.400000 83.365000 70.200000 84.615000 ;
        RECT 57.600000 99.645000 59.400000 100.895000 ;
        RECT 57.600000 107.785000 59.400000 109.035000 ;
        RECT 46.800000 107.785000 48.600000 109.035000 ;
        RECT 46.800000 99.645000 48.600000 100.895000 ;
        RECT 68.400000 107.785000 70.200000 109.035000 ;
        RECT 68.400000 99.645000 70.200000 100.895000 ;
        RECT 14.400000 132.205000 16.200000 133.455000 ;
        RECT 14.400000 124.065000 16.200000 125.315000 ;
        RECT 4.160000 124.065000 6.160000 125.315000 ;
        RECT 4.160000 132.205000 6.160000 133.455000 ;
        RECT 25.200000 132.205000 27.000000 133.455000 ;
        RECT 25.200000 124.065000 27.000000 125.315000 ;
        RECT 36.000000 124.065000 37.800000 125.315000 ;
        RECT 36.000000 132.205000 37.800000 133.455000 ;
        RECT 14.400000 148.485000 16.200000 149.735000 ;
        RECT 14.400000 140.345000 16.200000 141.595000 ;
        RECT 4.160000 140.345000 6.160000 141.595000 ;
        RECT 4.160000 148.485000 6.160000 149.735000 ;
        RECT 25.200000 140.345000 27.000000 141.595000 ;
        RECT 25.200000 148.485000 27.000000 149.735000 ;
        RECT 36.000000 140.345000 37.800000 141.595000 ;
        RECT 36.000000 148.485000 37.800000 149.735000 ;
        RECT 57.600000 124.065000 59.400000 125.315000 ;
        RECT 57.600000 132.205000 59.400000 133.455000 ;
        RECT 46.800000 132.205000 48.600000 133.455000 ;
        RECT 46.800000 124.065000 48.600000 125.315000 ;
        RECT 68.400000 132.205000 70.200000 133.455000 ;
        RECT 68.400000 124.065000 70.200000 125.315000 ;
        RECT 57.600000 140.345000 59.400000 141.595000 ;
        RECT 57.600000 148.485000 59.400000 149.735000 ;
        RECT 46.800000 148.485000 48.600000 149.735000 ;
        RECT 46.800000 140.345000 48.600000 141.595000 ;
        RECT 68.400000 148.485000 70.200000 149.735000 ;
        RECT 68.400000 140.345000 70.200000 141.595000 ;
        RECT 144.000000 115.925000 145.800000 117.175000 ;
        RECT 133.200000 115.925000 135.000000 117.175000 ;
        RECT 122.400000 115.925000 124.200000 117.175000 ;
        RECT 111.600000 115.925000 113.400000 117.175000 ;
        RECT 100.800000 115.925000 102.600000 117.175000 ;
        RECT 90.000000 115.925000 91.800000 117.175000 ;
        RECT 79.200000 115.925000 81.000000 117.175000 ;
        RECT 90.000000 91.505000 91.800000 92.755000 ;
        RECT 90.000000 83.365000 91.800000 84.615000 ;
        RECT 79.200000 83.365000 81.000000 84.615000 ;
        RECT 79.200000 91.505000 81.000000 92.755000 ;
        RECT 111.600000 91.505000 113.400000 92.755000 ;
        RECT 111.600000 83.365000 113.400000 84.615000 ;
        RECT 100.800000 91.505000 102.600000 92.755000 ;
        RECT 100.800000 83.365000 102.600000 84.615000 ;
        RECT 90.000000 107.785000 91.800000 109.035000 ;
        RECT 90.000000 99.645000 91.800000 100.895000 ;
        RECT 79.200000 107.785000 81.000000 109.035000 ;
        RECT 79.200000 99.645000 81.000000 100.895000 ;
        RECT 100.800000 107.785000 102.600000 109.035000 ;
        RECT 100.800000 99.645000 102.600000 100.895000 ;
        RECT 111.600000 99.645000 113.400000 100.895000 ;
        RECT 111.600000 107.785000 113.400000 109.035000 ;
        RECT 122.400000 83.365000 124.200000 84.615000 ;
        RECT 133.200000 83.365000 135.000000 84.615000 ;
        RECT 122.400000 91.505000 124.200000 92.755000 ;
        RECT 133.200000 91.505000 135.000000 92.755000 ;
        RECT 144.000000 91.505000 145.800000 92.755000 ;
        RECT 144.000000 83.365000 145.800000 84.615000 ;
        RECT 133.200000 107.785000 135.000000 109.035000 ;
        RECT 133.200000 99.645000 135.000000 100.895000 ;
        RECT 122.400000 107.785000 124.200000 109.035000 ;
        RECT 122.400000 99.645000 124.200000 100.895000 ;
        RECT 144.000000 107.785000 145.800000 109.035000 ;
        RECT 144.000000 99.645000 145.800000 100.895000 ;
        RECT 90.000000 132.205000 91.800000 133.455000 ;
        RECT 90.000000 124.065000 91.800000 125.315000 ;
        RECT 79.200000 124.065000 81.000000 125.315000 ;
        RECT 79.200000 132.205000 81.000000 133.455000 ;
        RECT 111.600000 132.205000 113.400000 133.455000 ;
        RECT 111.600000 124.065000 113.400000 125.315000 ;
        RECT 100.800000 132.205000 102.600000 133.455000 ;
        RECT 100.800000 124.065000 102.600000 125.315000 ;
        RECT 90.000000 148.485000 91.800000 149.735000 ;
        RECT 90.000000 140.345000 91.800000 141.595000 ;
        RECT 79.200000 148.485000 81.000000 149.735000 ;
        RECT 79.200000 140.345000 81.000000 141.595000 ;
        RECT 100.800000 148.485000 102.600000 149.735000 ;
        RECT 100.800000 140.345000 102.600000 141.595000 ;
        RECT 111.600000 140.345000 113.400000 141.595000 ;
        RECT 111.600000 148.485000 113.400000 149.735000 ;
        RECT 133.200000 132.205000 135.000000 133.455000 ;
        RECT 133.200000 124.065000 135.000000 125.315000 ;
        RECT 122.400000 132.205000 124.200000 133.455000 ;
        RECT 122.400000 124.065000 124.200000 125.315000 ;
        RECT 144.000000 132.205000 145.800000 133.455000 ;
        RECT 144.000000 124.065000 145.800000 125.315000 ;
        RECT 133.200000 148.485000 135.000000 149.735000 ;
        RECT 133.200000 140.345000 135.000000 141.595000 ;
        RECT 122.400000 148.485000 124.200000 149.735000 ;
        RECT 122.400000 140.345000 124.200000 141.595000 ;
        RECT 144.000000 148.485000 145.800000 149.735000 ;
        RECT 144.000000 140.345000 145.800000 141.595000 ;
        RECT 165.600000 75.225000 167.400000 76.475000 ;
        RECT 176.400000 75.225000 178.200000 76.475000 ;
        RECT 187.200000 75.225000 189.000000 76.475000 ;
        RECT 208.800000 75.225000 210.600000 76.475000 ;
        RECT 198.000000 75.225000 199.800000 76.475000 ;
        RECT 230.400000 75.225000 232.200000 76.475000 ;
        RECT 219.600000 75.225000 221.400000 76.475000 ;
        RECT 304.880000 18.245000 306.880000 19.495000 ;
        RECT 304.880000 10.615000 306.880000 11.355000 ;
        RECT 304.880000 26.385000 306.880000 27.635000 ;
        RECT 304.880000 34.525000 306.880000 35.775000 ;
        RECT 252.000000 75.225000 253.800000 76.475000 ;
        RECT 241.200000 75.225000 243.000000 76.475000 ;
        RECT 262.800000 75.225000 264.600000 76.475000 ;
        RECT 304.880000 42.665000 306.880000 43.915000 ;
        RECT 304.880000 50.805000 306.880000 52.055000 ;
        RECT 273.600000 75.225000 275.400000 76.475000 ;
        RECT 284.400000 75.225000 286.200000 76.475000 ;
        RECT 304.880000 75.225000 306.880000 76.475000 ;
        RECT 304.880000 67.085000 306.880000 68.335000 ;
        RECT 304.880000 58.945000 306.880000 60.195000 ;
        RECT 295.200000 75.225000 297.000000 76.475000 ;
        RECT 230.400000 115.925000 232.200000 117.175000 ;
        RECT 219.600000 115.925000 221.400000 117.175000 ;
        RECT 208.800000 115.925000 210.600000 117.175000 ;
        RECT 198.000000 115.925000 199.800000 117.175000 ;
        RECT 187.200000 115.925000 189.000000 117.175000 ;
        RECT 176.400000 115.925000 178.200000 117.175000 ;
        RECT 165.600000 115.925000 167.400000 117.175000 ;
        RECT 165.600000 83.365000 167.400000 84.615000 ;
        RECT 165.600000 91.505000 167.400000 92.755000 ;
        RECT 187.200000 91.505000 189.000000 92.755000 ;
        RECT 187.200000 83.365000 189.000000 84.615000 ;
        RECT 176.400000 91.505000 178.200000 92.755000 ;
        RECT 176.400000 83.365000 178.200000 84.615000 ;
        RECT 165.600000 107.785000 167.400000 109.035000 ;
        RECT 165.600000 99.645000 167.400000 100.895000 ;
        RECT 187.200000 107.785000 189.000000 109.035000 ;
        RECT 187.200000 99.645000 189.000000 100.895000 ;
        RECT 176.400000 107.785000 178.200000 109.035000 ;
        RECT 176.400000 99.645000 178.200000 100.895000 ;
        RECT 208.800000 91.505000 210.600000 92.755000 ;
        RECT 208.800000 83.365000 210.600000 84.615000 ;
        RECT 198.000000 91.505000 199.800000 92.755000 ;
        RECT 198.000000 83.365000 199.800000 84.615000 ;
        RECT 219.600000 83.365000 221.400000 84.615000 ;
        RECT 230.400000 83.365000 232.200000 84.615000 ;
        RECT 219.600000 91.505000 221.400000 92.755000 ;
        RECT 230.400000 91.505000 232.200000 92.755000 ;
        RECT 208.800000 107.785000 210.600000 109.035000 ;
        RECT 208.800000 99.645000 210.600000 100.895000 ;
        RECT 198.000000 107.785000 199.800000 109.035000 ;
        RECT 198.000000 99.645000 199.800000 100.895000 ;
        RECT 219.600000 107.785000 221.400000 109.035000 ;
        RECT 219.600000 99.645000 221.400000 100.895000 ;
        RECT 230.400000 99.645000 232.200000 100.895000 ;
        RECT 230.400000 107.785000 232.200000 109.035000 ;
        RECT 165.600000 124.065000 167.400000 125.315000 ;
        RECT 165.600000 132.205000 167.400000 133.455000 ;
        RECT 187.200000 132.205000 189.000000 133.455000 ;
        RECT 187.200000 124.065000 189.000000 125.315000 ;
        RECT 176.400000 132.205000 178.200000 133.455000 ;
        RECT 176.400000 124.065000 178.200000 125.315000 ;
        RECT 165.600000 148.485000 167.400000 149.735000 ;
        RECT 165.600000 140.345000 167.400000 141.595000 ;
        RECT 187.200000 148.485000 189.000000 149.735000 ;
        RECT 187.200000 140.345000 189.000000 141.595000 ;
        RECT 176.400000 148.485000 178.200000 149.735000 ;
        RECT 176.400000 140.345000 178.200000 141.595000 ;
        RECT 208.800000 132.205000 210.600000 133.455000 ;
        RECT 208.800000 124.065000 210.600000 125.315000 ;
        RECT 198.000000 132.205000 199.800000 133.455000 ;
        RECT 198.000000 124.065000 199.800000 125.315000 ;
        RECT 230.400000 132.205000 232.200000 133.455000 ;
        RECT 230.400000 124.065000 232.200000 125.315000 ;
        RECT 219.600000 132.205000 221.400000 133.455000 ;
        RECT 219.600000 124.065000 221.400000 125.315000 ;
        RECT 208.800000 148.485000 210.600000 149.735000 ;
        RECT 208.800000 140.345000 210.600000 141.595000 ;
        RECT 198.000000 148.485000 199.800000 149.735000 ;
        RECT 198.000000 140.345000 199.800000 141.595000 ;
        RECT 219.600000 148.485000 221.400000 149.735000 ;
        RECT 219.600000 140.345000 221.400000 141.595000 ;
        RECT 230.400000 140.345000 232.200000 141.595000 ;
        RECT 230.400000 148.485000 232.200000 149.735000 ;
        RECT 295.200000 115.925000 297.000000 117.175000 ;
        RECT 284.400000 115.925000 286.200000 117.175000 ;
        RECT 273.600000 115.925000 275.400000 117.175000 ;
        RECT 262.800000 115.925000 264.600000 117.175000 ;
        RECT 252.000000 115.925000 253.800000 117.175000 ;
        RECT 241.200000 115.925000 243.000000 117.175000 ;
        RECT 304.880000 115.925000 306.880000 117.175000 ;
        RECT 252.000000 83.365000 253.800000 84.615000 ;
        RECT 252.000000 91.505000 253.800000 92.755000 ;
        RECT 241.200000 91.505000 243.000000 92.755000 ;
        RECT 241.200000 83.365000 243.000000 84.615000 ;
        RECT 262.800000 91.505000 264.600000 92.755000 ;
        RECT 262.800000 83.365000 264.600000 84.615000 ;
        RECT 252.000000 99.645000 253.800000 100.895000 ;
        RECT 252.000000 107.785000 253.800000 109.035000 ;
        RECT 241.200000 107.785000 243.000000 109.035000 ;
        RECT 241.200000 99.645000 243.000000 100.895000 ;
        RECT 262.800000 107.785000 264.600000 109.035000 ;
        RECT 262.800000 99.645000 264.600000 100.895000 ;
        RECT 284.400000 91.505000 286.200000 92.755000 ;
        RECT 284.400000 83.365000 286.200000 84.615000 ;
        RECT 273.600000 91.505000 275.400000 92.755000 ;
        RECT 273.600000 83.365000 275.400000 84.615000 ;
        RECT 304.880000 91.505000 306.880000 92.755000 ;
        RECT 304.880000 83.365000 306.880000 84.615000 ;
        RECT 295.200000 83.365000 297.000000 84.615000 ;
        RECT 295.200000 91.505000 297.000000 92.755000 ;
        RECT 273.600000 107.785000 275.400000 109.035000 ;
        RECT 273.600000 99.645000 275.400000 100.895000 ;
        RECT 284.400000 99.645000 286.200000 100.895000 ;
        RECT 284.400000 107.785000 286.200000 109.035000 ;
        RECT 304.880000 107.785000 306.880000 109.035000 ;
        RECT 304.880000 99.645000 306.880000 100.895000 ;
        RECT 295.200000 99.645000 297.000000 100.895000 ;
        RECT 295.200000 107.785000 297.000000 109.035000 ;
        RECT 252.000000 124.065000 253.800000 125.315000 ;
        RECT 252.000000 132.205000 253.800000 133.455000 ;
        RECT 241.200000 132.205000 243.000000 133.455000 ;
        RECT 241.200000 124.065000 243.000000 125.315000 ;
        RECT 262.800000 132.205000 264.600000 133.455000 ;
        RECT 262.800000 124.065000 264.600000 125.315000 ;
        RECT 252.000000 140.345000 253.800000 141.595000 ;
        RECT 252.000000 148.485000 253.800000 149.735000 ;
        RECT 241.200000 148.485000 243.000000 149.735000 ;
        RECT 241.200000 140.345000 243.000000 141.595000 ;
        RECT 262.800000 148.485000 264.600000 149.735000 ;
        RECT 262.800000 140.345000 264.600000 141.595000 ;
        RECT 284.400000 132.205000 286.200000 133.455000 ;
        RECT 284.400000 124.065000 286.200000 125.315000 ;
        RECT 273.600000 132.205000 275.400000 133.455000 ;
        RECT 273.600000 124.065000 275.400000 125.315000 ;
        RECT 304.880000 124.065000 306.880000 125.315000 ;
        RECT 304.880000 132.205000 306.880000 133.455000 ;
        RECT 295.200000 124.065000 297.000000 125.315000 ;
        RECT 295.200000 132.205000 297.000000 133.455000 ;
        RECT 273.600000 148.485000 275.400000 149.735000 ;
        RECT 273.600000 140.345000 275.400000 141.595000 ;
        RECT 284.400000 140.345000 286.200000 141.595000 ;
        RECT 284.400000 148.485000 286.200000 149.735000 ;
        RECT 304.880000 140.345000 306.880000 141.595000 ;
        RECT 304.880000 148.485000 306.880000 149.735000 ;
        RECT 295.200000 140.345000 297.000000 141.595000 ;
        RECT 295.200000 148.485000 297.000000 149.735000 ;
        RECT 154.800000 156.625000 156.600000 157.875000 ;
        RECT 154.800000 164.765000 156.600000 166.015000 ;
        RECT 154.800000 172.905000 156.600000 174.155000 ;
        RECT 154.800000 181.045000 156.600000 182.295000 ;
        RECT 154.800000 189.185000 156.600000 190.435000 ;
        RECT 154.800000 213.605000 156.600000 214.855000 ;
        RECT 154.800000 197.325000 156.600000 198.575000 ;
        RECT 154.800000 205.465000 156.600000 206.715000 ;
        RECT 154.800000 221.745000 156.600000 222.995000 ;
        RECT 154.800000 229.885000 156.600000 231.135000 ;
        RECT 154.800000 238.025000 156.600000 239.275000 ;
        RECT 154.800000 246.165000 156.600000 247.415000 ;
        RECT 154.800000 254.305000 156.600000 255.555000 ;
        RECT 154.800000 262.445000 156.600000 263.695000 ;
        RECT 154.800000 270.585000 156.600000 271.835000 ;
        RECT 154.800000 278.725000 156.600000 279.975000 ;
        RECT 154.800000 286.865000 156.600000 288.115000 ;
        RECT 154.800000 295.005000 156.600000 296.255000 ;
        RECT 4.160000 164.765000 6.160000 166.015000 ;
        RECT 14.400000 164.765000 16.200000 166.015000 ;
        RECT 4.160000 156.625000 6.160000 157.875000 ;
        RECT 14.400000 156.625000 16.200000 157.875000 ;
        RECT 14.400000 172.905000 16.200000 174.155000 ;
        RECT 4.160000 172.905000 6.160000 174.155000 ;
        RECT 25.200000 164.765000 27.000000 166.015000 ;
        RECT 36.000000 164.765000 37.800000 166.015000 ;
        RECT 36.000000 156.625000 37.800000 157.875000 ;
        RECT 25.200000 156.625000 27.000000 157.875000 ;
        RECT 36.000000 172.905000 37.800000 174.155000 ;
        RECT 25.200000 172.905000 27.000000 174.155000 ;
        RECT 14.400000 181.045000 16.200000 182.295000 ;
        RECT 4.160000 181.045000 6.160000 182.295000 ;
        RECT 14.400000 189.185000 16.200000 190.435000 ;
        RECT 4.160000 189.185000 6.160000 190.435000 ;
        RECT 36.000000 181.045000 37.800000 182.295000 ;
        RECT 25.200000 181.045000 27.000000 182.295000 ;
        RECT 36.000000 189.185000 37.800000 190.435000 ;
        RECT 25.200000 189.185000 27.000000 190.435000 ;
        RECT 57.600000 156.625000 59.400000 157.875000 ;
        RECT 57.600000 164.765000 59.400000 166.015000 ;
        RECT 57.600000 172.905000 59.400000 174.155000 ;
        RECT 46.800000 172.905000 48.600000 174.155000 ;
        RECT 46.800000 164.765000 48.600000 166.015000 ;
        RECT 46.800000 156.625000 48.600000 157.875000 ;
        RECT 68.400000 172.905000 70.200000 174.155000 ;
        RECT 68.400000 164.765000 70.200000 166.015000 ;
        RECT 68.400000 156.625000 70.200000 157.875000 ;
        RECT 57.600000 181.045000 59.400000 182.295000 ;
        RECT 57.600000 189.185000 59.400000 190.435000 ;
        RECT 46.800000 189.185000 48.600000 190.435000 ;
        RECT 46.800000 181.045000 48.600000 182.295000 ;
        RECT 68.400000 189.185000 70.200000 190.435000 ;
        RECT 68.400000 181.045000 70.200000 182.295000 ;
        RECT 36.000000 213.605000 37.800000 214.855000 ;
        RECT 25.200000 213.605000 27.000000 214.855000 ;
        RECT 14.400000 213.605000 16.200000 214.855000 ;
        RECT 4.160000 213.605000 6.160000 214.855000 ;
        RECT 14.400000 197.325000 16.200000 198.575000 ;
        RECT 4.160000 205.465000 6.160000 206.715000 ;
        RECT 4.160000 197.325000 6.160000 198.575000 ;
        RECT 14.400000 205.465000 16.200000 206.715000 ;
        RECT 25.200000 197.325000 27.000000 198.575000 ;
        RECT 25.200000 205.465000 27.000000 206.715000 ;
        RECT 36.000000 197.325000 37.800000 198.575000 ;
        RECT 36.000000 205.465000 37.800000 206.715000 ;
        RECT 4.160000 229.885000 6.160000 231.135000 ;
        RECT 4.160000 221.745000 6.160000 222.995000 ;
        RECT 14.400000 221.745000 16.200000 222.995000 ;
        RECT 14.400000 229.885000 16.200000 231.135000 ;
        RECT 25.200000 221.745000 27.000000 222.995000 ;
        RECT 25.200000 229.885000 27.000000 231.135000 ;
        RECT 36.000000 221.745000 37.800000 222.995000 ;
        RECT 36.000000 229.885000 37.800000 231.135000 ;
        RECT 68.400000 213.605000 70.200000 214.855000 ;
        RECT 57.600000 213.605000 59.400000 214.855000 ;
        RECT 46.800000 213.605000 48.600000 214.855000 ;
        RECT 57.600000 197.325000 59.400000 198.575000 ;
        RECT 57.600000 205.465000 59.400000 206.715000 ;
        RECT 46.800000 205.465000 48.600000 206.715000 ;
        RECT 46.800000 197.325000 48.600000 198.575000 ;
        RECT 68.400000 205.465000 70.200000 206.715000 ;
        RECT 68.400000 197.325000 70.200000 198.575000 ;
        RECT 57.600000 221.745000 59.400000 222.995000 ;
        RECT 57.600000 229.885000 59.400000 231.135000 ;
        RECT 46.800000 229.885000 48.600000 231.135000 ;
        RECT 46.800000 221.745000 48.600000 222.995000 ;
        RECT 68.400000 229.885000 70.200000 231.135000 ;
        RECT 68.400000 221.745000 70.200000 222.995000 ;
        RECT 90.000000 172.905000 91.800000 174.155000 ;
        RECT 90.000000 164.765000 91.800000 166.015000 ;
        RECT 90.000000 156.625000 91.800000 157.875000 ;
        RECT 79.200000 172.905000 81.000000 174.155000 ;
        RECT 79.200000 164.765000 81.000000 166.015000 ;
        RECT 79.200000 156.625000 81.000000 157.875000 ;
        RECT 100.800000 156.625000 102.600000 157.875000 ;
        RECT 100.800000 164.765000 102.600000 166.015000 ;
        RECT 100.800000 172.905000 102.600000 174.155000 ;
        RECT 111.600000 156.625000 113.400000 157.875000 ;
        RECT 111.600000 164.765000 113.400000 166.015000 ;
        RECT 111.600000 172.905000 113.400000 174.155000 ;
        RECT 90.000000 189.185000 91.800000 190.435000 ;
        RECT 90.000000 181.045000 91.800000 182.295000 ;
        RECT 79.200000 189.185000 81.000000 190.435000 ;
        RECT 79.200000 181.045000 81.000000 182.295000 ;
        RECT 100.800000 181.045000 102.600000 182.295000 ;
        RECT 100.800000 189.185000 102.600000 190.435000 ;
        RECT 111.600000 181.045000 113.400000 182.295000 ;
        RECT 111.600000 189.185000 113.400000 190.435000 ;
        RECT 133.200000 164.765000 135.000000 166.015000 ;
        RECT 122.400000 164.765000 124.200000 166.015000 ;
        RECT 122.400000 156.625000 124.200000 157.875000 ;
        RECT 133.200000 156.625000 135.000000 157.875000 ;
        RECT 122.400000 172.905000 124.200000 174.155000 ;
        RECT 133.200000 172.905000 135.000000 174.155000 ;
        RECT 144.000000 172.905000 145.800000 174.155000 ;
        RECT 144.000000 164.765000 145.800000 166.015000 ;
        RECT 144.000000 156.625000 145.800000 157.875000 ;
        RECT 122.400000 181.045000 124.200000 182.295000 ;
        RECT 133.200000 181.045000 135.000000 182.295000 ;
        RECT 122.400000 189.185000 124.200000 190.435000 ;
        RECT 133.200000 189.185000 135.000000 190.435000 ;
        RECT 144.000000 189.185000 145.800000 190.435000 ;
        RECT 144.000000 181.045000 145.800000 182.295000 ;
        RECT 111.600000 213.605000 113.400000 214.855000 ;
        RECT 100.800000 213.605000 102.600000 214.855000 ;
        RECT 90.000000 213.605000 91.800000 214.855000 ;
        RECT 79.200000 213.605000 81.000000 214.855000 ;
        RECT 90.000000 205.465000 91.800000 206.715000 ;
        RECT 90.000000 197.325000 91.800000 198.575000 ;
        RECT 79.200000 205.465000 81.000000 206.715000 ;
        RECT 79.200000 197.325000 81.000000 198.575000 ;
        RECT 100.800000 197.325000 102.600000 198.575000 ;
        RECT 100.800000 205.465000 102.600000 206.715000 ;
        RECT 111.600000 197.325000 113.400000 198.575000 ;
        RECT 111.600000 205.465000 113.400000 206.715000 ;
        RECT 90.000000 229.885000 91.800000 231.135000 ;
        RECT 90.000000 221.745000 91.800000 222.995000 ;
        RECT 79.200000 229.885000 81.000000 231.135000 ;
        RECT 79.200000 221.745000 81.000000 222.995000 ;
        RECT 100.800000 221.745000 102.600000 222.995000 ;
        RECT 100.800000 229.885000 102.600000 231.135000 ;
        RECT 111.600000 221.745000 113.400000 222.995000 ;
        RECT 111.600000 229.885000 113.400000 231.135000 ;
        RECT 144.000000 213.605000 145.800000 214.855000 ;
        RECT 133.200000 213.605000 135.000000 214.855000 ;
        RECT 122.400000 213.605000 124.200000 214.855000 ;
        RECT 133.200000 205.465000 135.000000 206.715000 ;
        RECT 133.200000 197.325000 135.000000 198.575000 ;
        RECT 122.400000 205.465000 124.200000 206.715000 ;
        RECT 122.400000 197.325000 124.200000 198.575000 ;
        RECT 144.000000 205.465000 145.800000 206.715000 ;
        RECT 144.000000 197.325000 145.800000 198.575000 ;
        RECT 133.200000 229.885000 135.000000 231.135000 ;
        RECT 133.200000 221.745000 135.000000 222.995000 ;
        RECT 122.400000 229.885000 124.200000 231.135000 ;
        RECT 122.400000 221.745000 124.200000 222.995000 ;
        RECT 144.000000 229.885000 145.800000 231.135000 ;
        RECT 144.000000 221.745000 145.800000 222.995000 ;
        RECT 4.160000 238.025000 6.160000 239.275000 ;
        RECT 14.400000 238.025000 16.200000 239.275000 ;
        RECT 14.400000 246.165000 16.200000 247.415000 ;
        RECT 4.160000 246.165000 6.160000 247.415000 ;
        RECT 36.000000 238.025000 37.800000 239.275000 ;
        RECT 25.200000 238.025000 27.000000 239.275000 ;
        RECT 36.000000 246.165000 37.800000 247.415000 ;
        RECT 25.200000 246.165000 27.000000 247.415000 ;
        RECT 4.160000 262.445000 6.160000 263.695000 ;
        RECT 14.400000 262.445000 16.200000 263.695000 ;
        RECT 14.400000 254.305000 16.200000 255.555000 ;
        RECT 4.160000 254.305000 6.160000 255.555000 ;
        RECT 14.400000 270.585000 16.200000 271.835000 ;
        RECT 4.160000 270.585000 6.160000 271.835000 ;
        RECT 25.200000 262.445000 27.000000 263.695000 ;
        RECT 36.000000 262.445000 37.800000 263.695000 ;
        RECT 36.000000 254.305000 37.800000 255.555000 ;
        RECT 25.200000 254.305000 27.000000 255.555000 ;
        RECT 36.000000 270.585000 37.800000 271.835000 ;
        RECT 25.200000 270.585000 27.000000 271.835000 ;
        RECT 57.600000 238.025000 59.400000 239.275000 ;
        RECT 57.600000 246.165000 59.400000 247.415000 ;
        RECT 46.800000 246.165000 48.600000 247.415000 ;
        RECT 46.800000 238.025000 48.600000 239.275000 ;
        RECT 68.400000 246.165000 70.200000 247.415000 ;
        RECT 68.400000 238.025000 70.200000 239.275000 ;
        RECT 57.600000 254.305000 59.400000 255.555000 ;
        RECT 57.600000 262.445000 59.400000 263.695000 ;
        RECT 57.600000 270.585000 59.400000 271.835000 ;
        RECT 46.800000 270.585000 48.600000 271.835000 ;
        RECT 46.800000 262.445000 48.600000 263.695000 ;
        RECT 46.800000 254.305000 48.600000 255.555000 ;
        RECT 68.400000 270.585000 70.200000 271.835000 ;
        RECT 68.400000 262.445000 70.200000 263.695000 ;
        RECT 68.400000 254.305000 70.200000 255.555000 ;
        RECT 14.400000 286.865000 16.200000 288.115000 ;
        RECT 14.400000 278.725000 16.200000 279.975000 ;
        RECT 4.160000 278.725000 6.160000 279.975000 ;
        RECT 4.160000 286.865000 6.160000 288.115000 ;
        RECT 36.000000 286.865000 37.800000 288.115000 ;
        RECT 36.000000 278.725000 37.800000 279.975000 ;
        RECT 25.200000 286.865000 27.000000 288.115000 ;
        RECT 25.200000 278.725000 27.000000 279.975000 ;
        RECT 14.400000 295.005000 16.200000 296.255000 ;
        RECT 4.160000 295.005000 6.160000 296.255000 ;
        RECT 25.200000 295.005000 27.000000 296.255000 ;
        RECT 36.000000 295.005000 37.800000 296.255000 ;
        RECT 57.600000 278.725000 59.400000 279.975000 ;
        RECT 57.600000 286.865000 59.400000 288.115000 ;
        RECT 46.800000 286.865000 48.600000 288.115000 ;
        RECT 46.800000 278.725000 48.600000 279.975000 ;
        RECT 68.400000 286.865000 70.200000 288.115000 ;
        RECT 68.400000 278.725000 70.200000 279.975000 ;
        RECT 57.600000 295.005000 59.400000 296.255000 ;
        RECT 46.800000 295.005000 48.600000 296.255000 ;
        RECT 68.400000 295.005000 70.200000 296.255000 ;
        RECT 90.000000 246.165000 91.800000 247.415000 ;
        RECT 90.000000 238.025000 91.800000 239.275000 ;
        RECT 79.200000 246.165000 81.000000 247.415000 ;
        RECT 79.200000 238.025000 81.000000 239.275000 ;
        RECT 100.800000 238.025000 102.600000 239.275000 ;
        RECT 100.800000 246.165000 102.600000 247.415000 ;
        RECT 111.600000 238.025000 113.400000 239.275000 ;
        RECT 111.600000 246.165000 113.400000 247.415000 ;
        RECT 90.000000 270.585000 91.800000 271.835000 ;
        RECT 90.000000 262.445000 91.800000 263.695000 ;
        RECT 90.000000 254.305000 91.800000 255.555000 ;
        RECT 79.200000 270.585000 81.000000 271.835000 ;
        RECT 79.200000 262.445000 81.000000 263.695000 ;
        RECT 79.200000 254.305000 81.000000 255.555000 ;
        RECT 100.800000 254.305000 102.600000 255.555000 ;
        RECT 100.800000 262.445000 102.600000 263.695000 ;
        RECT 100.800000 270.585000 102.600000 271.835000 ;
        RECT 111.600000 254.305000 113.400000 255.555000 ;
        RECT 111.600000 262.445000 113.400000 263.695000 ;
        RECT 111.600000 270.585000 113.400000 271.835000 ;
        RECT 122.400000 238.025000 124.200000 239.275000 ;
        RECT 133.200000 238.025000 135.000000 239.275000 ;
        RECT 122.400000 246.165000 124.200000 247.415000 ;
        RECT 133.200000 246.165000 135.000000 247.415000 ;
        RECT 144.000000 246.165000 145.800000 247.415000 ;
        RECT 144.000000 238.025000 145.800000 239.275000 ;
        RECT 133.200000 262.445000 135.000000 263.695000 ;
        RECT 122.400000 262.445000 124.200000 263.695000 ;
        RECT 122.400000 254.305000 124.200000 255.555000 ;
        RECT 133.200000 254.305000 135.000000 255.555000 ;
        RECT 122.400000 270.585000 124.200000 271.835000 ;
        RECT 133.200000 270.585000 135.000000 271.835000 ;
        RECT 144.000000 270.585000 145.800000 271.835000 ;
        RECT 144.000000 262.445000 145.800000 263.695000 ;
        RECT 144.000000 254.305000 145.800000 255.555000 ;
        RECT 90.000000 286.865000 91.800000 288.115000 ;
        RECT 90.000000 278.725000 91.800000 279.975000 ;
        RECT 79.200000 278.725000 81.000000 279.975000 ;
        RECT 79.200000 286.865000 81.000000 288.115000 ;
        RECT 111.600000 286.865000 113.400000 288.115000 ;
        RECT 111.600000 278.725000 113.400000 279.975000 ;
        RECT 100.800000 286.865000 102.600000 288.115000 ;
        RECT 100.800000 278.725000 102.600000 279.975000 ;
        RECT 90.000000 295.005000 91.800000 296.255000 ;
        RECT 79.200000 295.005000 81.000000 296.255000 ;
        RECT 111.600000 295.005000 113.400000 296.255000 ;
        RECT 100.800000 295.005000 102.600000 296.255000 ;
        RECT 133.200000 286.865000 135.000000 288.115000 ;
        RECT 133.200000 278.725000 135.000000 279.975000 ;
        RECT 122.400000 286.865000 124.200000 288.115000 ;
        RECT 122.400000 278.725000 124.200000 279.975000 ;
        RECT 144.000000 286.865000 145.800000 288.115000 ;
        RECT 144.000000 278.725000 145.800000 279.975000 ;
        RECT 133.200000 295.005000 135.000000 296.255000 ;
        RECT 122.400000 295.005000 124.200000 296.255000 ;
        RECT 144.000000 295.005000 145.800000 296.255000 ;
        RECT 165.600000 172.905000 167.400000 174.155000 ;
        RECT 165.600000 164.765000 167.400000 166.015000 ;
        RECT 165.600000 156.625000 167.400000 157.875000 ;
        RECT 187.200000 172.905000 189.000000 174.155000 ;
        RECT 187.200000 164.765000 189.000000 166.015000 ;
        RECT 187.200000 156.625000 189.000000 157.875000 ;
        RECT 176.400000 172.905000 178.200000 174.155000 ;
        RECT 176.400000 164.765000 178.200000 166.015000 ;
        RECT 176.400000 156.625000 178.200000 157.875000 ;
        RECT 165.600000 189.185000 167.400000 190.435000 ;
        RECT 165.600000 181.045000 167.400000 182.295000 ;
        RECT 187.200000 189.185000 189.000000 190.435000 ;
        RECT 187.200000 181.045000 189.000000 182.295000 ;
        RECT 176.400000 189.185000 178.200000 190.435000 ;
        RECT 176.400000 181.045000 178.200000 182.295000 ;
        RECT 208.800000 172.905000 210.600000 174.155000 ;
        RECT 208.800000 164.765000 210.600000 166.015000 ;
        RECT 208.800000 156.625000 210.600000 157.875000 ;
        RECT 198.000000 172.905000 199.800000 174.155000 ;
        RECT 198.000000 164.765000 199.800000 166.015000 ;
        RECT 198.000000 156.625000 199.800000 157.875000 ;
        RECT 219.600000 164.765000 221.400000 166.015000 ;
        RECT 230.400000 164.765000 232.200000 166.015000 ;
        RECT 230.400000 156.625000 232.200000 157.875000 ;
        RECT 219.600000 156.625000 221.400000 157.875000 ;
        RECT 230.400000 172.905000 232.200000 174.155000 ;
        RECT 219.600000 172.905000 221.400000 174.155000 ;
        RECT 208.800000 189.185000 210.600000 190.435000 ;
        RECT 208.800000 181.045000 210.600000 182.295000 ;
        RECT 198.000000 189.185000 199.800000 190.435000 ;
        RECT 198.000000 181.045000 199.800000 182.295000 ;
        RECT 230.400000 181.045000 232.200000 182.295000 ;
        RECT 219.600000 181.045000 221.400000 182.295000 ;
        RECT 230.400000 189.185000 232.200000 190.435000 ;
        RECT 219.600000 189.185000 221.400000 190.435000 ;
        RECT 187.200000 213.605000 189.000000 214.855000 ;
        RECT 176.400000 213.605000 178.200000 214.855000 ;
        RECT 165.600000 213.605000 167.400000 214.855000 ;
        RECT 165.600000 205.465000 167.400000 206.715000 ;
        RECT 165.600000 197.325000 167.400000 198.575000 ;
        RECT 187.200000 205.465000 189.000000 206.715000 ;
        RECT 187.200000 197.325000 189.000000 198.575000 ;
        RECT 176.400000 205.465000 178.200000 206.715000 ;
        RECT 176.400000 197.325000 178.200000 198.575000 ;
        RECT 165.600000 229.885000 167.400000 231.135000 ;
        RECT 165.600000 221.745000 167.400000 222.995000 ;
        RECT 187.200000 229.885000 189.000000 231.135000 ;
        RECT 187.200000 221.745000 189.000000 222.995000 ;
        RECT 176.400000 229.885000 178.200000 231.135000 ;
        RECT 176.400000 221.745000 178.200000 222.995000 ;
        RECT 230.400000 213.605000 232.200000 214.855000 ;
        RECT 219.600000 213.605000 221.400000 214.855000 ;
        RECT 208.800000 213.605000 210.600000 214.855000 ;
        RECT 198.000000 213.605000 199.800000 214.855000 ;
        RECT 208.800000 205.465000 210.600000 206.715000 ;
        RECT 208.800000 197.325000 210.600000 198.575000 ;
        RECT 198.000000 205.465000 199.800000 206.715000 ;
        RECT 198.000000 197.325000 199.800000 198.575000 ;
        RECT 219.600000 197.325000 221.400000 198.575000 ;
        RECT 219.600000 205.465000 221.400000 206.715000 ;
        RECT 230.400000 197.325000 232.200000 198.575000 ;
        RECT 230.400000 205.465000 232.200000 206.715000 ;
        RECT 208.800000 229.885000 210.600000 231.135000 ;
        RECT 208.800000 221.745000 210.600000 222.995000 ;
        RECT 198.000000 229.885000 199.800000 231.135000 ;
        RECT 198.000000 221.745000 199.800000 222.995000 ;
        RECT 219.600000 221.745000 221.400000 222.995000 ;
        RECT 219.600000 229.885000 221.400000 231.135000 ;
        RECT 230.400000 221.745000 232.200000 222.995000 ;
        RECT 230.400000 229.885000 232.200000 231.135000 ;
        RECT 252.000000 156.625000 253.800000 157.875000 ;
        RECT 252.000000 164.765000 253.800000 166.015000 ;
        RECT 252.000000 172.905000 253.800000 174.155000 ;
        RECT 241.200000 172.905000 243.000000 174.155000 ;
        RECT 241.200000 164.765000 243.000000 166.015000 ;
        RECT 241.200000 156.625000 243.000000 157.875000 ;
        RECT 262.800000 172.905000 264.600000 174.155000 ;
        RECT 262.800000 164.765000 264.600000 166.015000 ;
        RECT 262.800000 156.625000 264.600000 157.875000 ;
        RECT 252.000000 181.045000 253.800000 182.295000 ;
        RECT 252.000000 189.185000 253.800000 190.435000 ;
        RECT 241.200000 189.185000 243.000000 190.435000 ;
        RECT 241.200000 181.045000 243.000000 182.295000 ;
        RECT 262.800000 189.185000 264.600000 190.435000 ;
        RECT 262.800000 181.045000 264.600000 182.295000 ;
        RECT 273.600000 156.625000 275.400000 157.875000 ;
        RECT 273.600000 164.765000 275.400000 166.015000 ;
        RECT 273.600000 172.905000 275.400000 174.155000 ;
        RECT 284.400000 156.625000 286.200000 157.875000 ;
        RECT 284.400000 164.765000 286.200000 166.015000 ;
        RECT 284.400000 172.905000 286.200000 174.155000 ;
        RECT 304.880000 172.905000 306.880000 174.155000 ;
        RECT 304.880000 164.765000 306.880000 166.015000 ;
        RECT 304.880000 156.625000 306.880000 157.875000 ;
        RECT 295.200000 156.625000 297.000000 157.875000 ;
        RECT 295.200000 164.765000 297.000000 166.015000 ;
        RECT 295.200000 172.905000 297.000000 174.155000 ;
        RECT 273.600000 181.045000 275.400000 182.295000 ;
        RECT 273.600000 189.185000 275.400000 190.435000 ;
        RECT 284.400000 181.045000 286.200000 182.295000 ;
        RECT 284.400000 189.185000 286.200000 190.435000 ;
        RECT 304.880000 189.185000 306.880000 190.435000 ;
        RECT 304.880000 181.045000 306.880000 182.295000 ;
        RECT 295.200000 181.045000 297.000000 182.295000 ;
        RECT 295.200000 189.185000 297.000000 190.435000 ;
        RECT 262.800000 213.605000 264.600000 214.855000 ;
        RECT 252.000000 213.605000 253.800000 214.855000 ;
        RECT 241.200000 213.605000 243.000000 214.855000 ;
        RECT 252.000000 197.325000 253.800000 198.575000 ;
        RECT 252.000000 205.465000 253.800000 206.715000 ;
        RECT 241.200000 205.465000 243.000000 206.715000 ;
        RECT 241.200000 197.325000 243.000000 198.575000 ;
        RECT 262.800000 205.465000 264.600000 206.715000 ;
        RECT 262.800000 197.325000 264.600000 198.575000 ;
        RECT 252.000000 221.745000 253.800000 222.995000 ;
        RECT 252.000000 229.885000 253.800000 231.135000 ;
        RECT 241.200000 229.885000 243.000000 231.135000 ;
        RECT 241.200000 221.745000 243.000000 222.995000 ;
        RECT 262.800000 229.885000 264.600000 231.135000 ;
        RECT 262.800000 221.745000 264.600000 222.995000 ;
        RECT 295.200000 213.605000 297.000000 214.855000 ;
        RECT 284.400000 213.605000 286.200000 214.855000 ;
        RECT 273.600000 213.605000 275.400000 214.855000 ;
        RECT 304.880000 213.605000 306.880000 214.855000 ;
        RECT 273.600000 197.325000 275.400000 198.575000 ;
        RECT 273.600000 205.465000 275.400000 206.715000 ;
        RECT 284.400000 197.325000 286.200000 198.575000 ;
        RECT 284.400000 205.465000 286.200000 206.715000 ;
        RECT 304.880000 205.465000 306.880000 206.715000 ;
        RECT 304.880000 197.325000 306.880000 198.575000 ;
        RECT 295.200000 197.325000 297.000000 198.575000 ;
        RECT 295.200000 205.465000 297.000000 206.715000 ;
        RECT 273.600000 221.745000 275.400000 222.995000 ;
        RECT 273.600000 229.885000 275.400000 231.135000 ;
        RECT 284.400000 221.745000 286.200000 222.995000 ;
        RECT 284.400000 229.885000 286.200000 231.135000 ;
        RECT 304.880000 229.885000 306.880000 231.135000 ;
        RECT 304.880000 221.745000 306.880000 222.995000 ;
        RECT 295.200000 221.745000 297.000000 222.995000 ;
        RECT 295.200000 229.885000 297.000000 231.135000 ;
        RECT 165.600000 246.165000 167.400000 247.415000 ;
        RECT 165.600000 238.025000 167.400000 239.275000 ;
        RECT 187.200000 246.165000 189.000000 247.415000 ;
        RECT 187.200000 238.025000 189.000000 239.275000 ;
        RECT 176.400000 246.165000 178.200000 247.415000 ;
        RECT 176.400000 238.025000 178.200000 239.275000 ;
        RECT 165.600000 270.585000 167.400000 271.835000 ;
        RECT 165.600000 262.445000 167.400000 263.695000 ;
        RECT 165.600000 254.305000 167.400000 255.555000 ;
        RECT 187.200000 270.585000 189.000000 271.835000 ;
        RECT 187.200000 262.445000 189.000000 263.695000 ;
        RECT 187.200000 254.305000 189.000000 255.555000 ;
        RECT 176.400000 270.585000 178.200000 271.835000 ;
        RECT 176.400000 262.445000 178.200000 263.695000 ;
        RECT 176.400000 254.305000 178.200000 255.555000 ;
        RECT 208.800000 246.165000 210.600000 247.415000 ;
        RECT 208.800000 238.025000 210.600000 239.275000 ;
        RECT 198.000000 246.165000 199.800000 247.415000 ;
        RECT 198.000000 238.025000 199.800000 239.275000 ;
        RECT 230.400000 238.025000 232.200000 239.275000 ;
        RECT 219.600000 238.025000 221.400000 239.275000 ;
        RECT 230.400000 246.165000 232.200000 247.415000 ;
        RECT 219.600000 246.165000 221.400000 247.415000 ;
        RECT 208.800000 270.585000 210.600000 271.835000 ;
        RECT 208.800000 262.445000 210.600000 263.695000 ;
        RECT 208.800000 254.305000 210.600000 255.555000 ;
        RECT 198.000000 270.585000 199.800000 271.835000 ;
        RECT 198.000000 262.445000 199.800000 263.695000 ;
        RECT 198.000000 254.305000 199.800000 255.555000 ;
        RECT 219.600000 262.445000 221.400000 263.695000 ;
        RECT 230.400000 262.445000 232.200000 263.695000 ;
        RECT 230.400000 254.305000 232.200000 255.555000 ;
        RECT 219.600000 254.305000 221.400000 255.555000 ;
        RECT 230.400000 270.585000 232.200000 271.835000 ;
        RECT 219.600000 270.585000 221.400000 271.835000 ;
        RECT 165.600000 278.725000 167.400000 279.975000 ;
        RECT 165.600000 286.865000 167.400000 288.115000 ;
        RECT 187.200000 286.865000 189.000000 288.115000 ;
        RECT 187.200000 278.725000 189.000000 279.975000 ;
        RECT 176.400000 286.865000 178.200000 288.115000 ;
        RECT 176.400000 278.725000 178.200000 279.975000 ;
        RECT 165.600000 295.005000 167.400000 296.255000 ;
        RECT 176.400000 295.005000 178.200000 296.255000 ;
        RECT 187.200000 295.005000 189.000000 296.255000 ;
        RECT 208.800000 286.865000 210.600000 288.115000 ;
        RECT 208.800000 278.725000 210.600000 279.975000 ;
        RECT 198.000000 286.865000 199.800000 288.115000 ;
        RECT 198.000000 278.725000 199.800000 279.975000 ;
        RECT 230.400000 286.865000 232.200000 288.115000 ;
        RECT 230.400000 278.725000 232.200000 279.975000 ;
        RECT 219.600000 286.865000 221.400000 288.115000 ;
        RECT 219.600000 278.725000 221.400000 279.975000 ;
        RECT 208.800000 295.005000 210.600000 296.255000 ;
        RECT 198.000000 295.005000 199.800000 296.255000 ;
        RECT 230.400000 295.005000 232.200000 296.255000 ;
        RECT 219.600000 295.005000 221.400000 296.255000 ;
        RECT 252.000000 238.025000 253.800000 239.275000 ;
        RECT 252.000000 246.165000 253.800000 247.415000 ;
        RECT 241.200000 246.165000 243.000000 247.415000 ;
        RECT 241.200000 238.025000 243.000000 239.275000 ;
        RECT 262.800000 246.165000 264.600000 247.415000 ;
        RECT 262.800000 238.025000 264.600000 239.275000 ;
        RECT 252.000000 254.305000 253.800000 255.555000 ;
        RECT 252.000000 262.445000 253.800000 263.695000 ;
        RECT 252.000000 270.585000 253.800000 271.835000 ;
        RECT 241.200000 270.585000 243.000000 271.835000 ;
        RECT 241.200000 262.445000 243.000000 263.695000 ;
        RECT 241.200000 254.305000 243.000000 255.555000 ;
        RECT 262.800000 270.585000 264.600000 271.835000 ;
        RECT 262.800000 262.445000 264.600000 263.695000 ;
        RECT 262.800000 254.305000 264.600000 255.555000 ;
        RECT 273.600000 238.025000 275.400000 239.275000 ;
        RECT 273.600000 246.165000 275.400000 247.415000 ;
        RECT 284.400000 238.025000 286.200000 239.275000 ;
        RECT 284.400000 246.165000 286.200000 247.415000 ;
        RECT 304.880000 238.025000 306.880000 239.275000 ;
        RECT 304.880000 246.165000 306.880000 247.415000 ;
        RECT 295.200000 238.025000 297.000000 239.275000 ;
        RECT 295.200000 246.165000 297.000000 247.415000 ;
        RECT 273.600000 254.305000 275.400000 255.555000 ;
        RECT 273.600000 262.445000 275.400000 263.695000 ;
        RECT 273.600000 270.585000 275.400000 271.835000 ;
        RECT 284.400000 254.305000 286.200000 255.555000 ;
        RECT 284.400000 262.445000 286.200000 263.695000 ;
        RECT 284.400000 270.585000 286.200000 271.835000 ;
        RECT 304.880000 254.305000 306.880000 255.555000 ;
        RECT 304.880000 262.445000 306.880000 263.695000 ;
        RECT 304.880000 270.585000 306.880000 271.835000 ;
        RECT 295.200000 254.305000 297.000000 255.555000 ;
        RECT 295.200000 262.445000 297.000000 263.695000 ;
        RECT 295.200000 270.585000 297.000000 271.835000 ;
        RECT 252.000000 278.725000 253.800000 279.975000 ;
        RECT 252.000000 286.865000 253.800000 288.115000 ;
        RECT 241.200000 286.865000 243.000000 288.115000 ;
        RECT 241.200000 278.725000 243.000000 279.975000 ;
        RECT 262.800000 286.865000 264.600000 288.115000 ;
        RECT 262.800000 278.725000 264.600000 279.975000 ;
        RECT 252.000000 295.005000 253.800000 296.255000 ;
        RECT 241.200000 295.005000 243.000000 296.255000 ;
        RECT 262.800000 295.005000 264.600000 296.255000 ;
        RECT 284.400000 286.865000 286.200000 288.115000 ;
        RECT 284.400000 278.725000 286.200000 279.975000 ;
        RECT 273.600000 286.865000 275.400000 288.115000 ;
        RECT 273.600000 278.725000 275.400000 279.975000 ;
        RECT 295.200000 286.865000 297.000000 288.115000 ;
        RECT 295.200000 278.725000 297.000000 279.975000 ;
        RECT 304.880000 278.725000 306.880000 279.975000 ;
        RECT 304.880000 286.865000 306.880000 288.115000 ;
        RECT 284.400000 295.005000 286.200000 296.255000 ;
        RECT 273.600000 295.005000 275.400000 296.255000 ;
        RECT 304.880000 295.005000 306.880000 296.255000 ;
        RECT 295.200000 295.005000 297.000000 296.255000 ;
      LAYER met3 ;
        RECT 0.000000 4.330000 311.040000 6.330000 ;
        RECT 0.000000 304.100000 311.040000 306.100000 ;
        RECT 154.800000 75.225000 156.600000 76.475000 ;
        RECT 154.800000 115.925000 156.600000 117.175000 ;
        RECT 154.800000 83.365000 156.600000 84.615000 ;
        RECT 154.800000 91.505000 156.600000 92.755000 ;
        RECT 154.800000 99.645000 156.600000 100.895000 ;
        RECT 154.800000 107.785000 156.600000 109.035000 ;
        RECT 154.800000 124.065000 156.600000 125.315000 ;
        RECT 154.800000 132.205000 156.600000 133.455000 ;
        RECT 154.800000 140.345000 156.600000 141.595000 ;
        RECT 154.800000 148.485000 156.600000 149.735000 ;
        RECT 4.160000 18.245000 6.160000 19.495000 ;
        RECT 4.160000 10.615000 6.160000 11.355000 ;
        RECT 4.160000 26.385000 6.160000 27.635000 ;
        RECT 4.160000 34.525000 6.160000 35.775000 ;
        RECT 4.160000 42.665000 6.160000 43.915000 ;
        RECT 4.160000 50.805000 6.160000 52.055000 ;
        RECT 4.160000 58.945000 6.160000 60.195000 ;
        RECT 4.160000 67.085000 6.160000 68.335000 ;
        RECT 4.160000 75.225000 6.160000 76.475000 ;
        RECT 14.400000 75.225000 16.200000 76.475000 ;
        RECT 36.000000 75.225000 37.800000 76.475000 ;
        RECT 25.200000 75.225000 27.000000 76.475000 ;
        RECT 57.600000 75.225000 59.400000 76.475000 ;
        RECT 46.800000 75.225000 48.600000 76.475000 ;
        RECT 68.400000 75.225000 70.200000 76.475000 ;
        RECT 90.000000 75.225000 91.800000 76.475000 ;
        RECT 79.200000 75.225000 81.000000 76.475000 ;
        RECT 111.600000 75.225000 113.400000 76.475000 ;
        RECT 100.800000 75.225000 102.600000 76.475000 ;
        RECT 133.200000 75.225000 135.000000 76.475000 ;
        RECT 122.400000 75.225000 124.200000 76.475000 ;
        RECT 144.000000 75.225000 145.800000 76.475000 ;
        RECT 68.400000 115.925000 70.200000 117.175000 ;
        RECT 57.600000 115.925000 59.400000 117.175000 ;
        RECT 46.800000 115.925000 48.600000 117.175000 ;
        RECT 36.000000 115.925000 37.800000 117.175000 ;
        RECT 25.200000 115.925000 27.000000 117.175000 ;
        RECT 14.400000 115.925000 16.200000 117.175000 ;
        RECT 4.160000 115.925000 6.160000 117.175000 ;
        RECT 14.400000 83.365000 16.200000 84.615000 ;
        RECT 4.160000 83.365000 6.160000 84.615000 ;
        RECT 14.400000 91.505000 16.200000 92.755000 ;
        RECT 4.160000 91.505000 6.160000 92.755000 ;
        RECT 36.000000 83.365000 37.800000 84.615000 ;
        RECT 25.200000 83.365000 27.000000 84.615000 ;
        RECT 36.000000 91.505000 37.800000 92.755000 ;
        RECT 25.200000 91.505000 27.000000 92.755000 ;
        RECT 14.400000 107.785000 16.200000 109.035000 ;
        RECT 4.160000 99.645000 6.160000 100.895000 ;
        RECT 4.160000 107.785000 6.160000 109.035000 ;
        RECT 14.400000 99.645000 16.200000 100.895000 ;
        RECT 25.200000 99.645000 27.000000 100.895000 ;
        RECT 25.200000 107.785000 27.000000 109.035000 ;
        RECT 36.000000 99.645000 37.800000 100.895000 ;
        RECT 36.000000 107.785000 37.800000 109.035000 ;
        RECT 57.600000 91.505000 59.400000 92.755000 ;
        RECT 57.600000 83.365000 59.400000 84.615000 ;
        RECT 46.800000 83.365000 48.600000 84.615000 ;
        RECT 46.800000 91.505000 48.600000 92.755000 ;
        RECT 68.400000 91.505000 70.200000 92.755000 ;
        RECT 68.400000 83.365000 70.200000 84.615000 ;
        RECT 57.600000 99.645000 59.400000 100.895000 ;
        RECT 57.600000 107.785000 59.400000 109.035000 ;
        RECT 46.800000 99.645000 48.600000 100.895000 ;
        RECT 46.800000 107.785000 48.600000 109.035000 ;
        RECT 68.400000 107.785000 70.200000 109.035000 ;
        RECT 68.400000 99.645000 70.200000 100.895000 ;
        RECT 4.160000 124.065000 6.160000 125.315000 ;
        RECT 4.160000 132.205000 6.160000 133.455000 ;
        RECT 14.400000 124.065000 16.200000 125.315000 ;
        RECT 14.400000 132.205000 16.200000 133.455000 ;
        RECT 25.200000 124.065000 27.000000 125.315000 ;
        RECT 25.200000 132.205000 27.000000 133.455000 ;
        RECT 36.000000 124.065000 37.800000 125.315000 ;
        RECT 36.000000 132.205000 37.800000 133.455000 ;
        RECT 4.160000 140.345000 6.160000 141.595000 ;
        RECT 4.160000 148.485000 6.160000 149.735000 ;
        RECT 14.400000 140.345000 16.200000 141.595000 ;
        RECT 14.400000 148.485000 16.200000 149.735000 ;
        RECT 25.200000 140.345000 27.000000 141.595000 ;
        RECT 25.200000 148.485000 27.000000 149.735000 ;
        RECT 36.000000 140.345000 37.800000 141.595000 ;
        RECT 36.000000 148.485000 37.800000 149.735000 ;
        RECT 57.600000 132.205000 59.400000 133.455000 ;
        RECT 57.600000 124.065000 59.400000 125.315000 ;
        RECT 46.800000 124.065000 48.600000 125.315000 ;
        RECT 46.800000 132.205000 48.600000 133.455000 ;
        RECT 68.400000 132.205000 70.200000 133.455000 ;
        RECT 68.400000 124.065000 70.200000 125.315000 ;
        RECT 57.600000 140.345000 59.400000 141.595000 ;
        RECT 57.600000 148.485000 59.400000 149.735000 ;
        RECT 46.800000 140.345000 48.600000 141.595000 ;
        RECT 46.800000 148.485000 48.600000 149.735000 ;
        RECT 68.400000 148.485000 70.200000 149.735000 ;
        RECT 68.400000 140.345000 70.200000 141.595000 ;
        RECT 144.000000 115.925000 145.800000 117.175000 ;
        RECT 133.200000 115.925000 135.000000 117.175000 ;
        RECT 122.400000 115.925000 124.200000 117.175000 ;
        RECT 111.600000 115.925000 113.400000 117.175000 ;
        RECT 100.800000 115.925000 102.600000 117.175000 ;
        RECT 90.000000 115.925000 91.800000 117.175000 ;
        RECT 79.200000 115.925000 81.000000 117.175000 ;
        RECT 90.000000 91.505000 91.800000 92.755000 ;
        RECT 90.000000 83.365000 91.800000 84.615000 ;
        RECT 79.200000 91.505000 81.000000 92.755000 ;
        RECT 79.200000 83.365000 81.000000 84.615000 ;
        RECT 111.600000 91.505000 113.400000 92.755000 ;
        RECT 111.600000 83.365000 113.400000 84.615000 ;
        RECT 100.800000 91.505000 102.600000 92.755000 ;
        RECT 100.800000 83.365000 102.600000 84.615000 ;
        RECT 90.000000 107.785000 91.800000 109.035000 ;
        RECT 90.000000 99.645000 91.800000 100.895000 ;
        RECT 79.200000 107.785000 81.000000 109.035000 ;
        RECT 79.200000 99.645000 81.000000 100.895000 ;
        RECT 111.600000 99.645000 113.400000 100.895000 ;
        RECT 100.800000 107.785000 102.600000 109.035000 ;
        RECT 100.800000 99.645000 102.600000 100.895000 ;
        RECT 111.600000 107.785000 113.400000 109.035000 ;
        RECT 133.200000 83.365000 135.000000 84.615000 ;
        RECT 122.400000 83.365000 124.200000 84.615000 ;
        RECT 133.200000 91.505000 135.000000 92.755000 ;
        RECT 122.400000 91.505000 124.200000 92.755000 ;
        RECT 144.000000 83.365000 145.800000 84.615000 ;
        RECT 144.000000 91.505000 145.800000 92.755000 ;
        RECT 122.400000 99.645000 124.200000 100.895000 ;
        RECT 122.400000 107.785000 124.200000 109.035000 ;
        RECT 133.200000 99.645000 135.000000 100.895000 ;
        RECT 133.200000 107.785000 135.000000 109.035000 ;
        RECT 144.000000 99.645000 145.800000 100.895000 ;
        RECT 144.000000 107.785000 145.800000 109.035000 ;
        RECT 90.000000 132.205000 91.800000 133.455000 ;
        RECT 90.000000 124.065000 91.800000 125.315000 ;
        RECT 79.200000 132.205000 81.000000 133.455000 ;
        RECT 79.200000 124.065000 81.000000 125.315000 ;
        RECT 100.800000 132.205000 102.600000 133.455000 ;
        RECT 100.800000 124.065000 102.600000 125.315000 ;
        RECT 111.600000 124.065000 113.400000 125.315000 ;
        RECT 111.600000 132.205000 113.400000 133.455000 ;
        RECT 90.000000 148.485000 91.800000 149.735000 ;
        RECT 90.000000 140.345000 91.800000 141.595000 ;
        RECT 79.200000 148.485000 81.000000 149.735000 ;
        RECT 79.200000 140.345000 81.000000 141.595000 ;
        RECT 100.800000 148.485000 102.600000 149.735000 ;
        RECT 100.800000 140.345000 102.600000 141.595000 ;
        RECT 111.600000 140.345000 113.400000 141.595000 ;
        RECT 111.600000 148.485000 113.400000 149.735000 ;
        RECT 122.400000 124.065000 124.200000 125.315000 ;
        RECT 122.400000 132.205000 124.200000 133.455000 ;
        RECT 133.200000 124.065000 135.000000 125.315000 ;
        RECT 133.200000 132.205000 135.000000 133.455000 ;
        RECT 144.000000 124.065000 145.800000 125.315000 ;
        RECT 144.000000 132.205000 145.800000 133.455000 ;
        RECT 122.400000 140.345000 124.200000 141.595000 ;
        RECT 122.400000 148.485000 124.200000 149.735000 ;
        RECT 133.200000 140.345000 135.000000 141.595000 ;
        RECT 133.200000 148.485000 135.000000 149.735000 ;
        RECT 144.000000 140.345000 145.800000 141.595000 ;
        RECT 144.000000 148.485000 145.800000 149.735000 ;
        RECT 176.400000 75.225000 178.200000 76.475000 ;
        RECT 165.600000 75.225000 167.400000 76.475000 ;
        RECT 187.200000 75.225000 189.000000 76.475000 ;
        RECT 208.800000 75.225000 210.600000 76.475000 ;
        RECT 198.000000 75.225000 199.800000 76.475000 ;
        RECT 230.400000 75.225000 232.200000 76.475000 ;
        RECT 219.600000 75.225000 221.400000 76.475000 ;
        RECT 304.880000 18.245000 306.880000 19.495000 ;
        RECT 304.880000 10.615000 306.880000 11.355000 ;
        RECT 304.880000 34.525000 306.880000 35.775000 ;
        RECT 304.880000 26.385000 306.880000 27.635000 ;
        RECT 252.000000 75.225000 253.800000 76.475000 ;
        RECT 241.200000 75.225000 243.000000 76.475000 ;
        RECT 262.800000 75.225000 264.600000 76.475000 ;
        RECT 304.880000 50.805000 306.880000 52.055000 ;
        RECT 304.880000 42.665000 306.880000 43.915000 ;
        RECT 273.600000 75.225000 275.400000 76.475000 ;
        RECT 284.400000 75.225000 286.200000 76.475000 ;
        RECT 304.880000 58.945000 306.880000 60.195000 ;
        RECT 304.880000 67.085000 306.880000 68.335000 ;
        RECT 304.880000 75.225000 306.880000 76.475000 ;
        RECT 295.200000 75.225000 297.000000 76.475000 ;
        RECT 230.400000 115.925000 232.200000 117.175000 ;
        RECT 219.600000 115.925000 221.400000 117.175000 ;
        RECT 208.800000 115.925000 210.600000 117.175000 ;
        RECT 198.000000 115.925000 199.800000 117.175000 ;
        RECT 187.200000 115.925000 189.000000 117.175000 ;
        RECT 176.400000 115.925000 178.200000 117.175000 ;
        RECT 165.600000 115.925000 167.400000 117.175000 ;
        RECT 165.600000 83.365000 167.400000 84.615000 ;
        RECT 165.600000 91.505000 167.400000 92.755000 ;
        RECT 187.200000 91.505000 189.000000 92.755000 ;
        RECT 187.200000 83.365000 189.000000 84.615000 ;
        RECT 176.400000 91.505000 178.200000 92.755000 ;
        RECT 176.400000 83.365000 178.200000 84.615000 ;
        RECT 165.600000 107.785000 167.400000 109.035000 ;
        RECT 165.600000 99.645000 167.400000 100.895000 ;
        RECT 187.200000 107.785000 189.000000 109.035000 ;
        RECT 187.200000 99.645000 189.000000 100.895000 ;
        RECT 176.400000 107.785000 178.200000 109.035000 ;
        RECT 176.400000 99.645000 178.200000 100.895000 ;
        RECT 198.000000 91.505000 199.800000 92.755000 ;
        RECT 198.000000 83.365000 199.800000 84.615000 ;
        RECT 208.800000 83.365000 210.600000 84.615000 ;
        RECT 208.800000 91.505000 210.600000 92.755000 ;
        RECT 230.400000 83.365000 232.200000 84.615000 ;
        RECT 219.600000 83.365000 221.400000 84.615000 ;
        RECT 230.400000 91.505000 232.200000 92.755000 ;
        RECT 219.600000 91.505000 221.400000 92.755000 ;
        RECT 198.000000 99.645000 199.800000 100.895000 ;
        RECT 198.000000 107.785000 199.800000 109.035000 ;
        RECT 208.800000 99.645000 210.600000 100.895000 ;
        RECT 208.800000 107.785000 210.600000 109.035000 ;
        RECT 219.600000 99.645000 221.400000 100.895000 ;
        RECT 219.600000 107.785000 221.400000 109.035000 ;
        RECT 230.400000 99.645000 232.200000 100.895000 ;
        RECT 230.400000 107.785000 232.200000 109.035000 ;
        RECT 165.600000 132.205000 167.400000 133.455000 ;
        RECT 165.600000 124.065000 167.400000 125.315000 ;
        RECT 187.200000 132.205000 189.000000 133.455000 ;
        RECT 187.200000 124.065000 189.000000 125.315000 ;
        RECT 176.400000 132.205000 178.200000 133.455000 ;
        RECT 176.400000 124.065000 178.200000 125.315000 ;
        RECT 165.600000 148.485000 167.400000 149.735000 ;
        RECT 165.600000 140.345000 167.400000 141.595000 ;
        RECT 187.200000 148.485000 189.000000 149.735000 ;
        RECT 187.200000 140.345000 189.000000 141.595000 ;
        RECT 176.400000 148.485000 178.200000 149.735000 ;
        RECT 176.400000 140.345000 178.200000 141.595000 ;
        RECT 198.000000 124.065000 199.800000 125.315000 ;
        RECT 198.000000 132.205000 199.800000 133.455000 ;
        RECT 208.800000 124.065000 210.600000 125.315000 ;
        RECT 208.800000 132.205000 210.600000 133.455000 ;
        RECT 219.600000 124.065000 221.400000 125.315000 ;
        RECT 219.600000 132.205000 221.400000 133.455000 ;
        RECT 230.400000 124.065000 232.200000 125.315000 ;
        RECT 230.400000 132.205000 232.200000 133.455000 ;
        RECT 198.000000 140.345000 199.800000 141.595000 ;
        RECT 198.000000 148.485000 199.800000 149.735000 ;
        RECT 208.800000 140.345000 210.600000 141.595000 ;
        RECT 208.800000 148.485000 210.600000 149.735000 ;
        RECT 219.600000 140.345000 221.400000 141.595000 ;
        RECT 219.600000 148.485000 221.400000 149.735000 ;
        RECT 230.400000 140.345000 232.200000 141.595000 ;
        RECT 230.400000 148.485000 232.200000 149.735000 ;
        RECT 295.200000 115.925000 297.000000 117.175000 ;
        RECT 284.400000 115.925000 286.200000 117.175000 ;
        RECT 273.600000 115.925000 275.400000 117.175000 ;
        RECT 262.800000 115.925000 264.600000 117.175000 ;
        RECT 252.000000 115.925000 253.800000 117.175000 ;
        RECT 241.200000 115.925000 243.000000 117.175000 ;
        RECT 304.880000 115.925000 306.880000 117.175000 ;
        RECT 252.000000 91.505000 253.800000 92.755000 ;
        RECT 252.000000 83.365000 253.800000 84.615000 ;
        RECT 241.200000 91.505000 243.000000 92.755000 ;
        RECT 241.200000 83.365000 243.000000 84.615000 ;
        RECT 262.800000 83.365000 264.600000 84.615000 ;
        RECT 262.800000 91.505000 264.600000 92.755000 ;
        RECT 252.000000 107.785000 253.800000 109.035000 ;
        RECT 252.000000 99.645000 253.800000 100.895000 ;
        RECT 241.200000 99.645000 243.000000 100.895000 ;
        RECT 241.200000 107.785000 243.000000 109.035000 ;
        RECT 262.800000 99.645000 264.600000 100.895000 ;
        RECT 262.800000 107.785000 264.600000 109.035000 ;
        RECT 273.600000 83.365000 275.400000 84.615000 ;
        RECT 273.600000 91.505000 275.400000 92.755000 ;
        RECT 284.400000 83.365000 286.200000 84.615000 ;
        RECT 284.400000 91.505000 286.200000 92.755000 ;
        RECT 295.200000 91.505000 297.000000 92.755000 ;
        RECT 295.200000 83.365000 297.000000 84.615000 ;
        RECT 304.880000 83.365000 306.880000 84.615000 ;
        RECT 304.880000 91.505000 306.880000 92.755000 ;
        RECT 284.400000 107.785000 286.200000 109.035000 ;
        RECT 284.400000 99.645000 286.200000 100.895000 ;
        RECT 273.600000 99.645000 275.400000 100.895000 ;
        RECT 273.600000 107.785000 275.400000 109.035000 ;
        RECT 295.200000 107.785000 297.000000 109.035000 ;
        RECT 295.200000 99.645000 297.000000 100.895000 ;
        RECT 304.880000 99.645000 306.880000 100.895000 ;
        RECT 304.880000 107.785000 306.880000 109.035000 ;
        RECT 252.000000 132.205000 253.800000 133.455000 ;
        RECT 252.000000 124.065000 253.800000 125.315000 ;
        RECT 241.200000 124.065000 243.000000 125.315000 ;
        RECT 241.200000 132.205000 243.000000 133.455000 ;
        RECT 262.800000 124.065000 264.600000 125.315000 ;
        RECT 262.800000 132.205000 264.600000 133.455000 ;
        RECT 252.000000 148.485000 253.800000 149.735000 ;
        RECT 252.000000 140.345000 253.800000 141.595000 ;
        RECT 241.200000 140.345000 243.000000 141.595000 ;
        RECT 241.200000 148.485000 243.000000 149.735000 ;
        RECT 262.800000 140.345000 264.600000 141.595000 ;
        RECT 262.800000 148.485000 264.600000 149.735000 ;
        RECT 273.600000 124.065000 275.400000 125.315000 ;
        RECT 273.600000 132.205000 275.400000 133.455000 ;
        RECT 284.400000 124.065000 286.200000 125.315000 ;
        RECT 284.400000 132.205000 286.200000 133.455000 ;
        RECT 295.200000 132.205000 297.000000 133.455000 ;
        RECT 295.200000 124.065000 297.000000 125.315000 ;
        RECT 304.880000 124.065000 306.880000 125.315000 ;
        RECT 304.880000 132.205000 306.880000 133.455000 ;
        RECT 284.400000 148.485000 286.200000 149.735000 ;
        RECT 284.400000 140.345000 286.200000 141.595000 ;
        RECT 273.600000 140.345000 275.400000 141.595000 ;
        RECT 273.600000 148.485000 275.400000 149.735000 ;
        RECT 295.200000 148.485000 297.000000 149.735000 ;
        RECT 295.200000 140.345000 297.000000 141.595000 ;
        RECT 304.880000 140.345000 306.880000 141.595000 ;
        RECT 304.880000 148.485000 306.880000 149.735000 ;
        RECT 154.800000 156.625000 156.600000 157.875000 ;
        RECT 154.800000 164.765000 156.600000 166.015000 ;
        RECT 154.800000 172.905000 156.600000 174.155000 ;
        RECT 154.800000 181.045000 156.600000 182.295000 ;
        RECT 154.800000 189.185000 156.600000 190.435000 ;
        RECT 154.800000 213.605000 156.600000 214.855000 ;
        RECT 154.800000 197.325000 156.600000 198.575000 ;
        RECT 154.800000 205.465000 156.600000 206.715000 ;
        RECT 154.800000 221.745000 156.600000 222.995000 ;
        RECT 154.800000 229.885000 156.600000 231.135000 ;
        RECT 154.800000 238.025000 156.600000 239.275000 ;
        RECT 154.800000 246.165000 156.600000 247.415000 ;
        RECT 154.800000 254.305000 156.600000 255.555000 ;
        RECT 154.800000 262.445000 156.600000 263.695000 ;
        RECT 154.800000 270.585000 156.600000 271.835000 ;
        RECT 154.800000 278.725000 156.600000 279.975000 ;
        RECT 154.800000 286.865000 156.600000 288.115000 ;
        RECT 154.800000 295.005000 156.600000 296.255000 ;
        RECT 4.160000 164.765000 6.160000 166.015000 ;
        RECT 14.400000 164.765000 16.200000 166.015000 ;
        RECT 4.160000 156.625000 6.160000 157.875000 ;
        RECT 14.400000 156.625000 16.200000 157.875000 ;
        RECT 14.400000 172.905000 16.200000 174.155000 ;
        RECT 4.160000 172.905000 6.160000 174.155000 ;
        RECT 25.200000 164.765000 27.000000 166.015000 ;
        RECT 36.000000 164.765000 37.800000 166.015000 ;
        RECT 36.000000 156.625000 37.800000 157.875000 ;
        RECT 25.200000 156.625000 27.000000 157.875000 ;
        RECT 36.000000 172.905000 37.800000 174.155000 ;
        RECT 25.200000 172.905000 27.000000 174.155000 ;
        RECT 14.400000 181.045000 16.200000 182.295000 ;
        RECT 4.160000 181.045000 6.160000 182.295000 ;
        RECT 14.400000 189.185000 16.200000 190.435000 ;
        RECT 4.160000 189.185000 6.160000 190.435000 ;
        RECT 36.000000 181.045000 37.800000 182.295000 ;
        RECT 25.200000 181.045000 27.000000 182.295000 ;
        RECT 36.000000 189.185000 37.800000 190.435000 ;
        RECT 25.200000 189.185000 27.000000 190.435000 ;
        RECT 57.600000 156.625000 59.400000 157.875000 ;
        RECT 57.600000 164.765000 59.400000 166.015000 ;
        RECT 57.600000 172.905000 59.400000 174.155000 ;
        RECT 46.800000 172.905000 48.600000 174.155000 ;
        RECT 46.800000 164.765000 48.600000 166.015000 ;
        RECT 46.800000 156.625000 48.600000 157.875000 ;
        RECT 68.400000 172.905000 70.200000 174.155000 ;
        RECT 68.400000 164.765000 70.200000 166.015000 ;
        RECT 68.400000 156.625000 70.200000 157.875000 ;
        RECT 57.600000 181.045000 59.400000 182.295000 ;
        RECT 57.600000 189.185000 59.400000 190.435000 ;
        RECT 46.800000 189.185000 48.600000 190.435000 ;
        RECT 46.800000 181.045000 48.600000 182.295000 ;
        RECT 68.400000 189.185000 70.200000 190.435000 ;
        RECT 68.400000 181.045000 70.200000 182.295000 ;
        RECT 4.160000 213.605000 6.160000 214.855000 ;
        RECT 14.400000 213.605000 16.200000 214.855000 ;
        RECT 25.200000 213.605000 27.000000 214.855000 ;
        RECT 36.000000 213.605000 37.800000 214.855000 ;
        RECT 4.160000 197.325000 6.160000 198.575000 ;
        RECT 4.160000 205.465000 6.160000 206.715000 ;
        RECT 14.400000 197.325000 16.200000 198.575000 ;
        RECT 14.400000 205.465000 16.200000 206.715000 ;
        RECT 25.200000 197.325000 27.000000 198.575000 ;
        RECT 25.200000 205.465000 27.000000 206.715000 ;
        RECT 36.000000 197.325000 37.800000 198.575000 ;
        RECT 36.000000 205.465000 37.800000 206.715000 ;
        RECT 4.160000 221.745000 6.160000 222.995000 ;
        RECT 4.160000 229.885000 6.160000 231.135000 ;
        RECT 14.400000 221.745000 16.200000 222.995000 ;
        RECT 14.400000 229.885000 16.200000 231.135000 ;
        RECT 25.200000 221.745000 27.000000 222.995000 ;
        RECT 25.200000 229.885000 27.000000 231.135000 ;
        RECT 36.000000 221.745000 37.800000 222.995000 ;
        RECT 36.000000 229.885000 37.800000 231.135000 ;
        RECT 68.400000 213.605000 70.200000 214.855000 ;
        RECT 57.600000 213.605000 59.400000 214.855000 ;
        RECT 46.800000 213.605000 48.600000 214.855000 ;
        RECT 57.600000 197.325000 59.400000 198.575000 ;
        RECT 57.600000 205.465000 59.400000 206.715000 ;
        RECT 46.800000 205.465000 48.600000 206.715000 ;
        RECT 46.800000 197.325000 48.600000 198.575000 ;
        RECT 68.400000 205.465000 70.200000 206.715000 ;
        RECT 68.400000 197.325000 70.200000 198.575000 ;
        RECT 57.600000 221.745000 59.400000 222.995000 ;
        RECT 57.600000 229.885000 59.400000 231.135000 ;
        RECT 46.800000 229.885000 48.600000 231.135000 ;
        RECT 46.800000 221.745000 48.600000 222.995000 ;
        RECT 68.400000 229.885000 70.200000 231.135000 ;
        RECT 68.400000 221.745000 70.200000 222.995000 ;
        RECT 90.000000 172.905000 91.800000 174.155000 ;
        RECT 90.000000 164.765000 91.800000 166.015000 ;
        RECT 90.000000 156.625000 91.800000 157.875000 ;
        RECT 79.200000 172.905000 81.000000 174.155000 ;
        RECT 79.200000 164.765000 81.000000 166.015000 ;
        RECT 79.200000 156.625000 81.000000 157.875000 ;
        RECT 100.800000 172.905000 102.600000 174.155000 ;
        RECT 100.800000 164.765000 102.600000 166.015000 ;
        RECT 100.800000 156.625000 102.600000 157.875000 ;
        RECT 111.600000 156.625000 113.400000 157.875000 ;
        RECT 111.600000 164.765000 113.400000 166.015000 ;
        RECT 111.600000 172.905000 113.400000 174.155000 ;
        RECT 90.000000 189.185000 91.800000 190.435000 ;
        RECT 90.000000 181.045000 91.800000 182.295000 ;
        RECT 79.200000 189.185000 81.000000 190.435000 ;
        RECT 79.200000 181.045000 81.000000 182.295000 ;
        RECT 100.800000 189.185000 102.600000 190.435000 ;
        RECT 100.800000 181.045000 102.600000 182.295000 ;
        RECT 111.600000 181.045000 113.400000 182.295000 ;
        RECT 111.600000 189.185000 113.400000 190.435000 ;
        RECT 122.400000 164.765000 124.200000 166.015000 ;
        RECT 133.200000 164.765000 135.000000 166.015000 ;
        RECT 133.200000 156.625000 135.000000 157.875000 ;
        RECT 122.400000 156.625000 124.200000 157.875000 ;
        RECT 133.200000 172.905000 135.000000 174.155000 ;
        RECT 122.400000 172.905000 124.200000 174.155000 ;
        RECT 144.000000 172.905000 145.800000 174.155000 ;
        RECT 144.000000 164.765000 145.800000 166.015000 ;
        RECT 144.000000 156.625000 145.800000 157.875000 ;
        RECT 133.200000 181.045000 135.000000 182.295000 ;
        RECT 122.400000 181.045000 124.200000 182.295000 ;
        RECT 133.200000 189.185000 135.000000 190.435000 ;
        RECT 122.400000 189.185000 124.200000 190.435000 ;
        RECT 144.000000 189.185000 145.800000 190.435000 ;
        RECT 144.000000 181.045000 145.800000 182.295000 ;
        RECT 100.800000 213.605000 102.600000 214.855000 ;
        RECT 90.000000 213.605000 91.800000 214.855000 ;
        RECT 79.200000 213.605000 81.000000 214.855000 ;
        RECT 111.600000 213.605000 113.400000 214.855000 ;
        RECT 90.000000 205.465000 91.800000 206.715000 ;
        RECT 90.000000 197.325000 91.800000 198.575000 ;
        RECT 79.200000 205.465000 81.000000 206.715000 ;
        RECT 79.200000 197.325000 81.000000 198.575000 ;
        RECT 100.800000 205.465000 102.600000 206.715000 ;
        RECT 100.800000 197.325000 102.600000 198.575000 ;
        RECT 111.600000 197.325000 113.400000 198.575000 ;
        RECT 111.600000 205.465000 113.400000 206.715000 ;
        RECT 90.000000 229.885000 91.800000 231.135000 ;
        RECT 90.000000 221.745000 91.800000 222.995000 ;
        RECT 79.200000 229.885000 81.000000 231.135000 ;
        RECT 79.200000 221.745000 81.000000 222.995000 ;
        RECT 100.800000 229.885000 102.600000 231.135000 ;
        RECT 100.800000 221.745000 102.600000 222.995000 ;
        RECT 111.600000 221.745000 113.400000 222.995000 ;
        RECT 111.600000 229.885000 113.400000 231.135000 ;
        RECT 144.000000 213.605000 145.800000 214.855000 ;
        RECT 122.400000 213.605000 124.200000 214.855000 ;
        RECT 133.200000 213.605000 135.000000 214.855000 ;
        RECT 122.400000 197.325000 124.200000 198.575000 ;
        RECT 122.400000 205.465000 124.200000 206.715000 ;
        RECT 133.200000 197.325000 135.000000 198.575000 ;
        RECT 133.200000 205.465000 135.000000 206.715000 ;
        RECT 144.000000 205.465000 145.800000 206.715000 ;
        RECT 144.000000 197.325000 145.800000 198.575000 ;
        RECT 122.400000 221.745000 124.200000 222.995000 ;
        RECT 122.400000 229.885000 124.200000 231.135000 ;
        RECT 133.200000 221.745000 135.000000 222.995000 ;
        RECT 133.200000 229.885000 135.000000 231.135000 ;
        RECT 144.000000 229.885000 145.800000 231.135000 ;
        RECT 144.000000 221.745000 145.800000 222.995000 ;
        RECT 14.400000 238.025000 16.200000 239.275000 ;
        RECT 4.160000 238.025000 6.160000 239.275000 ;
        RECT 14.400000 246.165000 16.200000 247.415000 ;
        RECT 4.160000 246.165000 6.160000 247.415000 ;
        RECT 36.000000 238.025000 37.800000 239.275000 ;
        RECT 25.200000 238.025000 27.000000 239.275000 ;
        RECT 36.000000 246.165000 37.800000 247.415000 ;
        RECT 25.200000 246.165000 27.000000 247.415000 ;
        RECT 4.160000 262.445000 6.160000 263.695000 ;
        RECT 14.400000 262.445000 16.200000 263.695000 ;
        RECT 14.400000 254.305000 16.200000 255.555000 ;
        RECT 4.160000 254.305000 6.160000 255.555000 ;
        RECT 14.400000 270.585000 16.200000 271.835000 ;
        RECT 4.160000 270.585000 6.160000 271.835000 ;
        RECT 25.200000 262.445000 27.000000 263.695000 ;
        RECT 36.000000 262.445000 37.800000 263.695000 ;
        RECT 36.000000 254.305000 37.800000 255.555000 ;
        RECT 25.200000 254.305000 27.000000 255.555000 ;
        RECT 36.000000 270.585000 37.800000 271.835000 ;
        RECT 25.200000 270.585000 27.000000 271.835000 ;
        RECT 57.600000 238.025000 59.400000 239.275000 ;
        RECT 57.600000 246.165000 59.400000 247.415000 ;
        RECT 46.800000 246.165000 48.600000 247.415000 ;
        RECT 46.800000 238.025000 48.600000 239.275000 ;
        RECT 68.400000 246.165000 70.200000 247.415000 ;
        RECT 68.400000 238.025000 70.200000 239.275000 ;
        RECT 57.600000 254.305000 59.400000 255.555000 ;
        RECT 57.600000 262.445000 59.400000 263.695000 ;
        RECT 57.600000 270.585000 59.400000 271.835000 ;
        RECT 46.800000 270.585000 48.600000 271.835000 ;
        RECT 46.800000 262.445000 48.600000 263.695000 ;
        RECT 46.800000 254.305000 48.600000 255.555000 ;
        RECT 68.400000 270.585000 70.200000 271.835000 ;
        RECT 68.400000 262.445000 70.200000 263.695000 ;
        RECT 68.400000 254.305000 70.200000 255.555000 ;
        RECT 4.160000 278.725000 6.160000 279.975000 ;
        RECT 4.160000 286.865000 6.160000 288.115000 ;
        RECT 14.400000 278.725000 16.200000 279.975000 ;
        RECT 14.400000 286.865000 16.200000 288.115000 ;
        RECT 25.200000 278.725000 27.000000 279.975000 ;
        RECT 25.200000 286.865000 27.000000 288.115000 ;
        RECT 36.000000 278.725000 37.800000 279.975000 ;
        RECT 36.000000 286.865000 37.800000 288.115000 ;
        RECT 4.160000 295.005000 6.160000 296.255000 ;
        RECT 14.400000 295.005000 16.200000 296.255000 ;
        RECT 25.200000 295.005000 27.000000 296.255000 ;
        RECT 36.000000 295.005000 37.800000 296.255000 ;
        RECT 57.600000 286.865000 59.400000 288.115000 ;
        RECT 57.600000 278.725000 59.400000 279.975000 ;
        RECT 46.800000 278.725000 48.600000 279.975000 ;
        RECT 46.800000 286.865000 48.600000 288.115000 ;
        RECT 68.400000 286.865000 70.200000 288.115000 ;
        RECT 68.400000 278.725000 70.200000 279.975000 ;
        RECT 57.600000 295.005000 59.400000 296.255000 ;
        RECT 46.800000 295.005000 48.600000 296.255000 ;
        RECT 68.400000 295.005000 70.200000 296.255000 ;
        RECT 90.000000 246.165000 91.800000 247.415000 ;
        RECT 90.000000 238.025000 91.800000 239.275000 ;
        RECT 79.200000 246.165000 81.000000 247.415000 ;
        RECT 79.200000 238.025000 81.000000 239.275000 ;
        RECT 100.800000 246.165000 102.600000 247.415000 ;
        RECT 100.800000 238.025000 102.600000 239.275000 ;
        RECT 111.600000 238.025000 113.400000 239.275000 ;
        RECT 111.600000 246.165000 113.400000 247.415000 ;
        RECT 90.000000 270.585000 91.800000 271.835000 ;
        RECT 90.000000 262.445000 91.800000 263.695000 ;
        RECT 90.000000 254.305000 91.800000 255.555000 ;
        RECT 79.200000 270.585000 81.000000 271.835000 ;
        RECT 79.200000 262.445000 81.000000 263.695000 ;
        RECT 79.200000 254.305000 81.000000 255.555000 ;
        RECT 100.800000 270.585000 102.600000 271.835000 ;
        RECT 100.800000 262.445000 102.600000 263.695000 ;
        RECT 100.800000 254.305000 102.600000 255.555000 ;
        RECT 111.600000 254.305000 113.400000 255.555000 ;
        RECT 111.600000 262.445000 113.400000 263.695000 ;
        RECT 111.600000 270.585000 113.400000 271.835000 ;
        RECT 133.200000 238.025000 135.000000 239.275000 ;
        RECT 122.400000 238.025000 124.200000 239.275000 ;
        RECT 133.200000 246.165000 135.000000 247.415000 ;
        RECT 122.400000 246.165000 124.200000 247.415000 ;
        RECT 144.000000 246.165000 145.800000 247.415000 ;
        RECT 144.000000 238.025000 145.800000 239.275000 ;
        RECT 122.400000 262.445000 124.200000 263.695000 ;
        RECT 133.200000 262.445000 135.000000 263.695000 ;
        RECT 133.200000 254.305000 135.000000 255.555000 ;
        RECT 122.400000 254.305000 124.200000 255.555000 ;
        RECT 133.200000 270.585000 135.000000 271.835000 ;
        RECT 122.400000 270.585000 124.200000 271.835000 ;
        RECT 144.000000 270.585000 145.800000 271.835000 ;
        RECT 144.000000 262.445000 145.800000 263.695000 ;
        RECT 144.000000 254.305000 145.800000 255.555000 ;
        RECT 90.000000 286.865000 91.800000 288.115000 ;
        RECT 90.000000 278.725000 91.800000 279.975000 ;
        RECT 79.200000 286.865000 81.000000 288.115000 ;
        RECT 79.200000 278.725000 81.000000 279.975000 ;
        RECT 100.800000 286.865000 102.600000 288.115000 ;
        RECT 100.800000 278.725000 102.600000 279.975000 ;
        RECT 111.600000 278.725000 113.400000 279.975000 ;
        RECT 111.600000 286.865000 113.400000 288.115000 ;
        RECT 90.000000 295.005000 91.800000 296.255000 ;
        RECT 79.200000 295.005000 81.000000 296.255000 ;
        RECT 100.800000 295.005000 102.600000 296.255000 ;
        RECT 111.600000 295.005000 113.400000 296.255000 ;
        RECT 122.400000 278.725000 124.200000 279.975000 ;
        RECT 122.400000 286.865000 124.200000 288.115000 ;
        RECT 133.200000 278.725000 135.000000 279.975000 ;
        RECT 133.200000 286.865000 135.000000 288.115000 ;
        RECT 144.000000 278.725000 145.800000 279.975000 ;
        RECT 144.000000 286.865000 145.800000 288.115000 ;
        RECT 122.400000 295.005000 124.200000 296.255000 ;
        RECT 133.200000 295.005000 135.000000 296.255000 ;
        RECT 144.000000 295.005000 145.800000 296.255000 ;
        RECT 165.600000 172.905000 167.400000 174.155000 ;
        RECT 165.600000 164.765000 167.400000 166.015000 ;
        RECT 165.600000 156.625000 167.400000 157.875000 ;
        RECT 187.200000 172.905000 189.000000 174.155000 ;
        RECT 187.200000 164.765000 189.000000 166.015000 ;
        RECT 187.200000 156.625000 189.000000 157.875000 ;
        RECT 176.400000 172.905000 178.200000 174.155000 ;
        RECT 176.400000 164.765000 178.200000 166.015000 ;
        RECT 176.400000 156.625000 178.200000 157.875000 ;
        RECT 165.600000 189.185000 167.400000 190.435000 ;
        RECT 165.600000 181.045000 167.400000 182.295000 ;
        RECT 187.200000 189.185000 189.000000 190.435000 ;
        RECT 187.200000 181.045000 189.000000 182.295000 ;
        RECT 176.400000 189.185000 178.200000 190.435000 ;
        RECT 176.400000 181.045000 178.200000 182.295000 ;
        RECT 198.000000 156.625000 199.800000 157.875000 ;
        RECT 198.000000 164.765000 199.800000 166.015000 ;
        RECT 198.000000 172.905000 199.800000 174.155000 ;
        RECT 208.800000 156.625000 210.600000 157.875000 ;
        RECT 208.800000 164.765000 210.600000 166.015000 ;
        RECT 208.800000 172.905000 210.600000 174.155000 ;
        RECT 230.400000 164.765000 232.200000 166.015000 ;
        RECT 219.600000 164.765000 221.400000 166.015000 ;
        RECT 219.600000 156.625000 221.400000 157.875000 ;
        RECT 230.400000 156.625000 232.200000 157.875000 ;
        RECT 219.600000 172.905000 221.400000 174.155000 ;
        RECT 230.400000 172.905000 232.200000 174.155000 ;
        RECT 198.000000 181.045000 199.800000 182.295000 ;
        RECT 198.000000 189.185000 199.800000 190.435000 ;
        RECT 208.800000 181.045000 210.600000 182.295000 ;
        RECT 208.800000 189.185000 210.600000 190.435000 ;
        RECT 219.600000 181.045000 221.400000 182.295000 ;
        RECT 230.400000 181.045000 232.200000 182.295000 ;
        RECT 219.600000 189.185000 221.400000 190.435000 ;
        RECT 230.400000 189.185000 232.200000 190.435000 ;
        RECT 187.200000 213.605000 189.000000 214.855000 ;
        RECT 176.400000 213.605000 178.200000 214.855000 ;
        RECT 165.600000 213.605000 167.400000 214.855000 ;
        RECT 165.600000 205.465000 167.400000 206.715000 ;
        RECT 165.600000 197.325000 167.400000 198.575000 ;
        RECT 187.200000 205.465000 189.000000 206.715000 ;
        RECT 187.200000 197.325000 189.000000 198.575000 ;
        RECT 176.400000 205.465000 178.200000 206.715000 ;
        RECT 176.400000 197.325000 178.200000 198.575000 ;
        RECT 165.600000 229.885000 167.400000 231.135000 ;
        RECT 165.600000 221.745000 167.400000 222.995000 ;
        RECT 187.200000 229.885000 189.000000 231.135000 ;
        RECT 187.200000 221.745000 189.000000 222.995000 ;
        RECT 176.400000 229.885000 178.200000 231.135000 ;
        RECT 176.400000 221.745000 178.200000 222.995000 ;
        RECT 230.400000 213.605000 232.200000 214.855000 ;
        RECT 198.000000 213.605000 199.800000 214.855000 ;
        RECT 208.800000 213.605000 210.600000 214.855000 ;
        RECT 219.600000 213.605000 221.400000 214.855000 ;
        RECT 198.000000 197.325000 199.800000 198.575000 ;
        RECT 198.000000 205.465000 199.800000 206.715000 ;
        RECT 208.800000 197.325000 210.600000 198.575000 ;
        RECT 208.800000 205.465000 210.600000 206.715000 ;
        RECT 230.400000 205.465000 232.200000 206.715000 ;
        RECT 230.400000 197.325000 232.200000 198.575000 ;
        RECT 219.600000 197.325000 221.400000 198.575000 ;
        RECT 219.600000 205.465000 221.400000 206.715000 ;
        RECT 198.000000 221.745000 199.800000 222.995000 ;
        RECT 198.000000 229.885000 199.800000 231.135000 ;
        RECT 208.800000 221.745000 210.600000 222.995000 ;
        RECT 208.800000 229.885000 210.600000 231.135000 ;
        RECT 230.400000 229.885000 232.200000 231.135000 ;
        RECT 230.400000 221.745000 232.200000 222.995000 ;
        RECT 219.600000 221.745000 221.400000 222.995000 ;
        RECT 219.600000 229.885000 221.400000 231.135000 ;
        RECT 252.000000 172.905000 253.800000 174.155000 ;
        RECT 252.000000 164.765000 253.800000 166.015000 ;
        RECT 252.000000 156.625000 253.800000 157.875000 ;
        RECT 241.200000 156.625000 243.000000 157.875000 ;
        RECT 241.200000 164.765000 243.000000 166.015000 ;
        RECT 241.200000 172.905000 243.000000 174.155000 ;
        RECT 262.800000 156.625000 264.600000 157.875000 ;
        RECT 262.800000 164.765000 264.600000 166.015000 ;
        RECT 262.800000 172.905000 264.600000 174.155000 ;
        RECT 252.000000 189.185000 253.800000 190.435000 ;
        RECT 252.000000 181.045000 253.800000 182.295000 ;
        RECT 241.200000 181.045000 243.000000 182.295000 ;
        RECT 241.200000 189.185000 243.000000 190.435000 ;
        RECT 262.800000 181.045000 264.600000 182.295000 ;
        RECT 262.800000 189.185000 264.600000 190.435000 ;
        RECT 284.400000 172.905000 286.200000 174.155000 ;
        RECT 284.400000 164.765000 286.200000 166.015000 ;
        RECT 284.400000 156.625000 286.200000 157.875000 ;
        RECT 273.600000 172.905000 275.400000 174.155000 ;
        RECT 273.600000 164.765000 275.400000 166.015000 ;
        RECT 273.600000 156.625000 275.400000 157.875000 ;
        RECT 295.200000 172.905000 297.000000 174.155000 ;
        RECT 295.200000 164.765000 297.000000 166.015000 ;
        RECT 295.200000 156.625000 297.000000 157.875000 ;
        RECT 304.880000 156.625000 306.880000 157.875000 ;
        RECT 304.880000 164.765000 306.880000 166.015000 ;
        RECT 304.880000 172.905000 306.880000 174.155000 ;
        RECT 284.400000 189.185000 286.200000 190.435000 ;
        RECT 284.400000 181.045000 286.200000 182.295000 ;
        RECT 273.600000 189.185000 275.400000 190.435000 ;
        RECT 273.600000 181.045000 275.400000 182.295000 ;
        RECT 295.200000 189.185000 297.000000 190.435000 ;
        RECT 295.200000 181.045000 297.000000 182.295000 ;
        RECT 304.880000 181.045000 306.880000 182.295000 ;
        RECT 304.880000 189.185000 306.880000 190.435000 ;
        RECT 241.200000 213.605000 243.000000 214.855000 ;
        RECT 252.000000 213.605000 253.800000 214.855000 ;
        RECT 262.800000 213.605000 264.600000 214.855000 ;
        RECT 252.000000 205.465000 253.800000 206.715000 ;
        RECT 252.000000 197.325000 253.800000 198.575000 ;
        RECT 241.200000 197.325000 243.000000 198.575000 ;
        RECT 241.200000 205.465000 243.000000 206.715000 ;
        RECT 262.800000 197.325000 264.600000 198.575000 ;
        RECT 262.800000 205.465000 264.600000 206.715000 ;
        RECT 252.000000 229.885000 253.800000 231.135000 ;
        RECT 252.000000 221.745000 253.800000 222.995000 ;
        RECT 241.200000 221.745000 243.000000 222.995000 ;
        RECT 241.200000 229.885000 243.000000 231.135000 ;
        RECT 262.800000 221.745000 264.600000 222.995000 ;
        RECT 262.800000 229.885000 264.600000 231.135000 ;
        RECT 295.200000 213.605000 297.000000 214.855000 ;
        RECT 284.400000 213.605000 286.200000 214.855000 ;
        RECT 273.600000 213.605000 275.400000 214.855000 ;
        RECT 304.880000 213.605000 306.880000 214.855000 ;
        RECT 284.400000 205.465000 286.200000 206.715000 ;
        RECT 284.400000 197.325000 286.200000 198.575000 ;
        RECT 273.600000 205.465000 275.400000 206.715000 ;
        RECT 273.600000 197.325000 275.400000 198.575000 ;
        RECT 295.200000 205.465000 297.000000 206.715000 ;
        RECT 295.200000 197.325000 297.000000 198.575000 ;
        RECT 304.880000 197.325000 306.880000 198.575000 ;
        RECT 304.880000 205.465000 306.880000 206.715000 ;
        RECT 284.400000 229.885000 286.200000 231.135000 ;
        RECT 284.400000 221.745000 286.200000 222.995000 ;
        RECT 273.600000 229.885000 275.400000 231.135000 ;
        RECT 273.600000 221.745000 275.400000 222.995000 ;
        RECT 295.200000 229.885000 297.000000 231.135000 ;
        RECT 295.200000 221.745000 297.000000 222.995000 ;
        RECT 304.880000 221.745000 306.880000 222.995000 ;
        RECT 304.880000 229.885000 306.880000 231.135000 ;
        RECT 165.600000 246.165000 167.400000 247.415000 ;
        RECT 165.600000 238.025000 167.400000 239.275000 ;
        RECT 187.200000 246.165000 189.000000 247.415000 ;
        RECT 187.200000 238.025000 189.000000 239.275000 ;
        RECT 176.400000 246.165000 178.200000 247.415000 ;
        RECT 176.400000 238.025000 178.200000 239.275000 ;
        RECT 165.600000 270.585000 167.400000 271.835000 ;
        RECT 165.600000 262.445000 167.400000 263.695000 ;
        RECT 165.600000 254.305000 167.400000 255.555000 ;
        RECT 187.200000 270.585000 189.000000 271.835000 ;
        RECT 187.200000 262.445000 189.000000 263.695000 ;
        RECT 187.200000 254.305000 189.000000 255.555000 ;
        RECT 176.400000 270.585000 178.200000 271.835000 ;
        RECT 176.400000 262.445000 178.200000 263.695000 ;
        RECT 176.400000 254.305000 178.200000 255.555000 ;
        RECT 198.000000 238.025000 199.800000 239.275000 ;
        RECT 198.000000 246.165000 199.800000 247.415000 ;
        RECT 208.800000 238.025000 210.600000 239.275000 ;
        RECT 208.800000 246.165000 210.600000 247.415000 ;
        RECT 219.600000 238.025000 221.400000 239.275000 ;
        RECT 230.400000 238.025000 232.200000 239.275000 ;
        RECT 219.600000 246.165000 221.400000 247.415000 ;
        RECT 230.400000 246.165000 232.200000 247.415000 ;
        RECT 198.000000 254.305000 199.800000 255.555000 ;
        RECT 198.000000 262.445000 199.800000 263.695000 ;
        RECT 198.000000 270.585000 199.800000 271.835000 ;
        RECT 208.800000 254.305000 210.600000 255.555000 ;
        RECT 208.800000 262.445000 210.600000 263.695000 ;
        RECT 208.800000 270.585000 210.600000 271.835000 ;
        RECT 230.400000 262.445000 232.200000 263.695000 ;
        RECT 219.600000 262.445000 221.400000 263.695000 ;
        RECT 219.600000 254.305000 221.400000 255.555000 ;
        RECT 230.400000 254.305000 232.200000 255.555000 ;
        RECT 219.600000 270.585000 221.400000 271.835000 ;
        RECT 230.400000 270.585000 232.200000 271.835000 ;
        RECT 165.600000 286.865000 167.400000 288.115000 ;
        RECT 165.600000 278.725000 167.400000 279.975000 ;
        RECT 187.200000 286.865000 189.000000 288.115000 ;
        RECT 187.200000 278.725000 189.000000 279.975000 ;
        RECT 176.400000 286.865000 178.200000 288.115000 ;
        RECT 176.400000 278.725000 178.200000 279.975000 ;
        RECT 187.200000 295.005000 189.000000 296.255000 ;
        RECT 165.600000 295.005000 167.400000 296.255000 ;
        RECT 176.400000 295.005000 178.200000 296.255000 ;
        RECT 198.000000 278.725000 199.800000 279.975000 ;
        RECT 198.000000 286.865000 199.800000 288.115000 ;
        RECT 208.800000 278.725000 210.600000 279.975000 ;
        RECT 208.800000 286.865000 210.600000 288.115000 ;
        RECT 219.600000 278.725000 221.400000 279.975000 ;
        RECT 219.600000 286.865000 221.400000 288.115000 ;
        RECT 230.400000 278.725000 232.200000 279.975000 ;
        RECT 230.400000 286.865000 232.200000 288.115000 ;
        RECT 198.000000 295.005000 199.800000 296.255000 ;
        RECT 208.800000 295.005000 210.600000 296.255000 ;
        RECT 219.600000 295.005000 221.400000 296.255000 ;
        RECT 230.400000 295.005000 232.200000 296.255000 ;
        RECT 252.000000 246.165000 253.800000 247.415000 ;
        RECT 252.000000 238.025000 253.800000 239.275000 ;
        RECT 241.200000 238.025000 243.000000 239.275000 ;
        RECT 241.200000 246.165000 243.000000 247.415000 ;
        RECT 262.800000 238.025000 264.600000 239.275000 ;
        RECT 262.800000 246.165000 264.600000 247.415000 ;
        RECT 252.000000 270.585000 253.800000 271.835000 ;
        RECT 252.000000 262.445000 253.800000 263.695000 ;
        RECT 252.000000 254.305000 253.800000 255.555000 ;
        RECT 241.200000 254.305000 243.000000 255.555000 ;
        RECT 241.200000 262.445000 243.000000 263.695000 ;
        RECT 241.200000 270.585000 243.000000 271.835000 ;
        RECT 262.800000 254.305000 264.600000 255.555000 ;
        RECT 262.800000 262.445000 264.600000 263.695000 ;
        RECT 262.800000 270.585000 264.600000 271.835000 ;
        RECT 284.400000 246.165000 286.200000 247.415000 ;
        RECT 284.400000 238.025000 286.200000 239.275000 ;
        RECT 273.600000 246.165000 275.400000 247.415000 ;
        RECT 273.600000 238.025000 275.400000 239.275000 ;
        RECT 295.200000 246.165000 297.000000 247.415000 ;
        RECT 295.200000 238.025000 297.000000 239.275000 ;
        RECT 304.880000 238.025000 306.880000 239.275000 ;
        RECT 304.880000 246.165000 306.880000 247.415000 ;
        RECT 284.400000 270.585000 286.200000 271.835000 ;
        RECT 284.400000 262.445000 286.200000 263.695000 ;
        RECT 284.400000 254.305000 286.200000 255.555000 ;
        RECT 273.600000 270.585000 275.400000 271.835000 ;
        RECT 273.600000 262.445000 275.400000 263.695000 ;
        RECT 273.600000 254.305000 275.400000 255.555000 ;
        RECT 295.200000 270.585000 297.000000 271.835000 ;
        RECT 295.200000 262.445000 297.000000 263.695000 ;
        RECT 295.200000 254.305000 297.000000 255.555000 ;
        RECT 304.880000 254.305000 306.880000 255.555000 ;
        RECT 304.880000 262.445000 306.880000 263.695000 ;
        RECT 304.880000 270.585000 306.880000 271.835000 ;
        RECT 252.000000 286.865000 253.800000 288.115000 ;
        RECT 252.000000 278.725000 253.800000 279.975000 ;
        RECT 241.200000 278.725000 243.000000 279.975000 ;
        RECT 241.200000 286.865000 243.000000 288.115000 ;
        RECT 262.800000 278.725000 264.600000 279.975000 ;
        RECT 262.800000 286.865000 264.600000 288.115000 ;
        RECT 252.000000 295.005000 253.800000 296.255000 ;
        RECT 241.200000 295.005000 243.000000 296.255000 ;
        RECT 262.800000 295.005000 264.600000 296.255000 ;
        RECT 273.600000 278.725000 275.400000 279.975000 ;
        RECT 273.600000 286.865000 275.400000 288.115000 ;
        RECT 284.400000 278.725000 286.200000 279.975000 ;
        RECT 284.400000 286.865000 286.200000 288.115000 ;
        RECT 295.200000 286.865000 297.000000 288.115000 ;
        RECT 295.200000 278.725000 297.000000 279.975000 ;
        RECT 304.880000 278.725000 306.880000 279.975000 ;
        RECT 304.880000 286.865000 306.880000 288.115000 ;
        RECT 284.400000 295.005000 286.200000 296.255000 ;
        RECT 273.600000 295.005000 275.400000 296.255000 ;
        RECT 295.200000 295.005000 297.000000 296.255000 ;
        RECT 304.880000 295.005000 306.880000 296.255000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VREG
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 154.800000 0.000000 156.800000 3.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.400000 0.000000 16.200000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.200000 0.000000 27.000000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.000000 0.000000 37.800000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.800000 0.000000 48.600000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.600000 0.000000 59.400000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.400000 0.000000 70.200000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.200000 0.000000 81.000000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 90.000000 0.000000 91.800000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.800000 0.000000 102.600000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 111.600000 0.000000 113.400000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.400000 0.000000 124.200000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 133.200000 0.000000 135.000000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.000000 0.000000 145.800000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.800000 0.000000 156.600000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.600000 0.000000 167.400000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 176.400000 0.000000 178.200000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 187.200000 0.000000 189.000000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 198.000000 0.000000 199.800000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.800000 0.000000 210.600000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.600000 0.000000 221.400000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 230.400000 0.000000 232.200000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 241.200000 0.000000 243.000000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 252.000000 0.000000 253.800000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 262.800000 0.000000 264.600000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 273.600000 0.000000 275.400000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.400000 0.000000 286.200000 1.800000 ;
    END
    PORT
      LAYER met4 ;
        RECT 295.200000 0.000000 297.000000 1.800000 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.040000 307.300000 311.040000 309.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 307.300000 2.000000 309.300000 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.040000 1.130000 311.040000 3.130000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 1.130000 2.000000 3.130000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.080000 309.540000 310.080000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.080000 0.000000 310.080000 2.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.960000 309.540000 2.960000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.960000 0.000000 2.960000 2.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 0.000000 1.130000 311.040000 3.130000 ;
        RECT 0.000000 307.300000 311.040000 309.300000 ;
    END
# end of P/G power stripe data as pin

  END VREG
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 309.040000 300.900000 311.040000 302.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 300.900000 2.000000 302.900000 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.040000 7.530000 311.040000 9.530000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000000 7.530000 2.000000 9.530000 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.680000 309.540000 303.680000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.680000 0.000000 303.680000 2.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.360000 309.540000 9.360000 311.540000 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.360000 0.000000 9.360000 2.000000 ;
    END

# P/G power stripe data as pin
    PORT
      LAYER met2 ;
        RECT 7.360000 38.595000 9.360000 39.845000 ;
        RECT 10.560000 38.595000 12.360000 39.845000 ;
        RECT 21.360000 38.595000 23.160000 39.845000 ;
        RECT 32.160000 38.595000 33.960000 39.845000 ;
        RECT 42.960000 38.595000 44.760000 39.845000 ;
        RECT 53.760000 38.595000 55.560000 39.845000 ;
        RECT 64.560000 38.595000 66.360000 39.845000 ;
        RECT 75.360000 38.595000 77.160000 39.845000 ;
        RECT 32.160000 14.175000 33.960000 15.425000 ;
        RECT 21.360000 14.175000 23.160000 15.425000 ;
        RECT 10.560000 14.175000 12.360000 15.425000 ;
        RECT 7.360000 14.175000 9.360000 15.425000 ;
        RECT 7.360000 22.315000 9.360000 23.565000 ;
        RECT 7.360000 30.455000 9.360000 31.705000 ;
        RECT 10.560000 22.315000 12.360000 23.565000 ;
        RECT 10.560000 30.455000 12.360000 31.705000 ;
        RECT 21.360000 22.315000 23.160000 23.565000 ;
        RECT 21.360000 30.455000 23.160000 31.705000 ;
        RECT 32.160000 22.315000 33.960000 23.565000 ;
        RECT 32.160000 30.455000 33.960000 31.705000 ;
        RECT 42.960000 14.175000 44.760000 15.425000 ;
        RECT 53.760000 14.175000 55.560000 15.425000 ;
        RECT 64.560000 14.175000 66.360000 15.425000 ;
        RECT 75.360000 14.175000 77.160000 15.425000 ;
        RECT 75.360000 30.455000 77.160000 31.705000 ;
        RECT 42.960000 22.315000 44.760000 23.565000 ;
        RECT 42.960000 30.455000 44.760000 31.705000 ;
        RECT 53.760000 22.315000 55.560000 23.565000 ;
        RECT 53.760000 30.455000 55.560000 31.705000 ;
        RECT 64.560000 22.315000 66.360000 23.565000 ;
        RECT 64.560000 30.455000 66.360000 31.705000 ;
        RECT 75.360000 22.315000 77.160000 23.565000 ;
        RECT 7.360000 54.875000 9.360000 56.125000 ;
        RECT 7.360000 46.735000 9.360000 47.985000 ;
        RECT 10.560000 46.735000 12.360000 47.985000 ;
        RECT 10.560000 54.875000 12.360000 56.125000 ;
        RECT 21.360000 46.735000 23.160000 47.985000 ;
        RECT 21.360000 54.875000 23.160000 56.125000 ;
        RECT 32.160000 46.735000 33.960000 47.985000 ;
        RECT 32.160000 54.875000 33.960000 56.125000 ;
        RECT 10.560000 71.155000 12.360000 72.405000 ;
        RECT 10.560000 63.015000 12.360000 64.265000 ;
        RECT 7.360000 63.015000 9.360000 64.265000 ;
        RECT 7.360000 71.155000 9.360000 72.405000 ;
        RECT 32.160000 71.155000 33.960000 72.405000 ;
        RECT 32.160000 63.015000 33.960000 64.265000 ;
        RECT 21.360000 71.155000 23.160000 72.405000 ;
        RECT 21.360000 63.015000 23.160000 64.265000 ;
        RECT 75.360000 54.875000 77.160000 56.125000 ;
        RECT 75.360000 46.735000 77.160000 47.985000 ;
        RECT 64.560000 54.875000 66.360000 56.125000 ;
        RECT 64.560000 46.735000 66.360000 47.985000 ;
        RECT 53.760000 54.875000 55.560000 56.125000 ;
        RECT 42.960000 46.735000 44.760000 47.985000 ;
        RECT 42.960000 54.875000 44.760000 56.125000 ;
        RECT 53.760000 46.735000 55.560000 47.985000 ;
        RECT 42.960000 71.155000 44.760000 72.405000 ;
        RECT 42.960000 63.015000 44.760000 64.265000 ;
        RECT 53.760000 63.015000 55.560000 64.265000 ;
        RECT 53.760000 71.155000 55.560000 72.405000 ;
        RECT 64.560000 63.015000 66.360000 64.265000 ;
        RECT 64.560000 71.155000 66.360000 72.405000 ;
        RECT 75.360000 63.015000 77.160000 64.265000 ;
        RECT 75.360000 71.155000 77.160000 72.405000 ;
        RECT 150.960000 38.595000 152.760000 39.845000 ;
        RECT 140.160000 38.595000 141.960000 39.845000 ;
        RECT 129.360000 38.595000 131.160000 39.845000 ;
        RECT 118.560000 38.595000 120.360000 39.845000 ;
        RECT 107.760000 38.595000 109.560000 39.845000 ;
        RECT 96.960000 38.595000 98.760000 39.845000 ;
        RECT 86.160000 38.595000 87.960000 39.845000 ;
        RECT 86.160000 14.175000 87.960000 15.425000 ;
        RECT 96.960000 14.175000 98.760000 15.425000 ;
        RECT 107.760000 14.175000 109.560000 15.425000 ;
        RECT 86.160000 22.315000 87.960000 23.565000 ;
        RECT 86.160000 30.455000 87.960000 31.705000 ;
        RECT 96.960000 22.315000 98.760000 23.565000 ;
        RECT 96.960000 30.455000 98.760000 31.705000 ;
        RECT 107.760000 22.315000 109.560000 23.565000 ;
        RECT 107.760000 30.455000 109.560000 31.705000 ;
        RECT 118.560000 14.175000 120.360000 15.425000 ;
        RECT 129.360000 14.175000 131.160000 15.425000 ;
        RECT 140.160000 14.175000 141.960000 15.425000 ;
        RECT 150.960000 14.175000 152.760000 15.425000 ;
        RECT 150.960000 30.455000 152.760000 31.705000 ;
        RECT 118.560000 22.315000 120.360000 23.565000 ;
        RECT 118.560000 30.455000 120.360000 31.705000 ;
        RECT 129.360000 22.315000 131.160000 23.565000 ;
        RECT 129.360000 30.455000 131.160000 31.705000 ;
        RECT 140.160000 22.315000 141.960000 23.565000 ;
        RECT 140.160000 30.455000 141.960000 31.705000 ;
        RECT 150.960000 22.315000 152.760000 23.565000 ;
        RECT 107.760000 54.875000 109.560000 56.125000 ;
        RECT 107.760000 46.735000 109.560000 47.985000 ;
        RECT 86.160000 46.735000 87.960000 47.985000 ;
        RECT 86.160000 54.875000 87.960000 56.125000 ;
        RECT 96.960000 46.735000 98.760000 47.985000 ;
        RECT 96.960000 54.875000 98.760000 56.125000 ;
        RECT 96.960000 71.155000 98.760000 72.405000 ;
        RECT 96.960000 63.015000 98.760000 64.265000 ;
        RECT 86.160000 71.155000 87.960000 72.405000 ;
        RECT 86.160000 63.015000 87.960000 64.265000 ;
        RECT 107.760000 63.015000 109.560000 64.265000 ;
        RECT 107.760000 71.155000 109.560000 72.405000 ;
        RECT 150.960000 54.875000 152.760000 56.125000 ;
        RECT 150.960000 46.735000 152.760000 47.985000 ;
        RECT 140.160000 54.875000 141.960000 56.125000 ;
        RECT 140.160000 46.735000 141.960000 47.985000 ;
        RECT 129.360000 54.875000 131.160000 56.125000 ;
        RECT 118.560000 46.735000 120.360000 47.985000 ;
        RECT 118.560000 54.875000 120.360000 56.125000 ;
        RECT 129.360000 46.735000 131.160000 47.985000 ;
        RECT 118.560000 71.155000 120.360000 72.405000 ;
        RECT 118.560000 63.015000 120.360000 64.265000 ;
        RECT 129.360000 63.015000 131.160000 64.265000 ;
        RECT 129.360000 71.155000 131.160000 72.405000 ;
        RECT 140.160000 63.015000 141.960000 64.265000 ;
        RECT 140.160000 71.155000 141.960000 72.405000 ;
        RECT 150.960000 63.015000 152.760000 64.265000 ;
        RECT 150.960000 71.155000 152.760000 72.405000 ;
        RECT 10.560000 87.435000 12.360000 88.685000 ;
        RECT 7.360000 87.435000 9.360000 88.685000 ;
        RECT 7.360000 79.295000 9.360000 80.545000 ;
        RECT 10.560000 79.295000 12.360000 80.545000 ;
        RECT 7.360000 95.575000 9.360000 96.825000 ;
        RECT 10.560000 95.575000 12.360000 96.825000 ;
        RECT 32.160000 87.435000 33.960000 88.685000 ;
        RECT 21.360000 87.435000 23.160000 88.685000 ;
        RECT 21.360000 79.295000 23.160000 80.545000 ;
        RECT 32.160000 79.295000 33.960000 80.545000 ;
        RECT 21.360000 95.575000 23.160000 96.825000 ;
        RECT 32.160000 95.575000 33.960000 96.825000 ;
        RECT 10.560000 111.855000 12.360000 113.105000 ;
        RECT 10.560000 103.715000 12.360000 104.965000 ;
        RECT 7.360000 103.715000 9.360000 104.965000 ;
        RECT 7.360000 111.855000 9.360000 113.105000 ;
        RECT 32.160000 111.855000 33.960000 113.105000 ;
        RECT 32.160000 103.715000 33.960000 104.965000 ;
        RECT 21.360000 111.855000 23.160000 113.105000 ;
        RECT 21.360000 103.715000 23.160000 104.965000 ;
        RECT 53.760000 95.575000 55.560000 96.825000 ;
        RECT 53.760000 87.435000 55.560000 88.685000 ;
        RECT 53.760000 79.295000 55.560000 80.545000 ;
        RECT 42.960000 95.575000 44.760000 96.825000 ;
        RECT 42.960000 87.435000 44.760000 88.685000 ;
        RECT 42.960000 79.295000 44.760000 80.545000 ;
        RECT 75.360000 95.575000 77.160000 96.825000 ;
        RECT 75.360000 87.435000 77.160000 88.685000 ;
        RECT 75.360000 79.295000 77.160000 80.545000 ;
        RECT 64.560000 95.575000 66.360000 96.825000 ;
        RECT 64.560000 87.435000 66.360000 88.685000 ;
        RECT 64.560000 79.295000 66.360000 80.545000 ;
        RECT 42.960000 103.715000 44.760000 104.965000 ;
        RECT 42.960000 111.855000 44.760000 113.105000 ;
        RECT 53.760000 103.715000 55.560000 104.965000 ;
        RECT 53.760000 111.855000 55.560000 113.105000 ;
        RECT 75.360000 111.855000 77.160000 113.105000 ;
        RECT 75.360000 103.715000 77.160000 104.965000 ;
        RECT 64.560000 111.855000 66.360000 113.105000 ;
        RECT 64.560000 103.715000 66.360000 104.965000 ;
        RECT 32.160000 136.275000 33.960000 137.525000 ;
        RECT 21.360000 136.275000 23.160000 137.525000 ;
        RECT 10.560000 136.275000 12.360000 137.525000 ;
        RECT 7.360000 136.275000 9.360000 137.525000 ;
        RECT 10.560000 128.135000 12.360000 129.385000 ;
        RECT 10.560000 119.995000 12.360000 121.245000 ;
        RECT 7.360000 119.995000 9.360000 121.245000 ;
        RECT 7.360000 128.135000 9.360000 129.385000 ;
        RECT 32.160000 128.135000 33.960000 129.385000 ;
        RECT 32.160000 119.995000 33.960000 121.245000 ;
        RECT 21.360000 128.135000 23.160000 129.385000 ;
        RECT 21.360000 119.995000 23.160000 121.245000 ;
        RECT 10.560000 152.555000 12.360000 153.805000 ;
        RECT 10.560000 144.415000 12.360000 145.665000 ;
        RECT 7.360000 144.415000 9.360000 145.665000 ;
        RECT 7.360000 152.555000 9.360000 153.805000 ;
        RECT 32.160000 152.555000 33.960000 153.805000 ;
        RECT 32.160000 144.415000 33.960000 145.665000 ;
        RECT 21.360000 152.555000 23.160000 153.805000 ;
        RECT 21.360000 144.415000 23.160000 145.665000 ;
        RECT 75.360000 136.275000 77.160000 137.525000 ;
        RECT 64.560000 136.275000 66.360000 137.525000 ;
        RECT 53.760000 136.275000 55.560000 137.525000 ;
        RECT 42.960000 136.275000 44.760000 137.525000 ;
        RECT 42.960000 119.995000 44.760000 121.245000 ;
        RECT 42.960000 128.135000 44.760000 129.385000 ;
        RECT 53.760000 119.995000 55.560000 121.245000 ;
        RECT 53.760000 128.135000 55.560000 129.385000 ;
        RECT 75.360000 128.135000 77.160000 129.385000 ;
        RECT 75.360000 119.995000 77.160000 121.245000 ;
        RECT 64.560000 128.135000 66.360000 129.385000 ;
        RECT 64.560000 119.995000 66.360000 121.245000 ;
        RECT 42.960000 144.415000 44.760000 145.665000 ;
        RECT 42.960000 152.555000 44.760000 153.805000 ;
        RECT 53.760000 144.415000 55.560000 145.665000 ;
        RECT 53.760000 152.555000 55.560000 153.805000 ;
        RECT 75.360000 152.555000 77.160000 153.805000 ;
        RECT 75.360000 144.415000 77.160000 145.665000 ;
        RECT 64.560000 152.555000 66.360000 153.805000 ;
        RECT 64.560000 144.415000 66.360000 145.665000 ;
        RECT 96.960000 95.575000 98.760000 96.825000 ;
        RECT 96.960000 87.435000 98.760000 88.685000 ;
        RECT 96.960000 79.295000 98.760000 80.545000 ;
        RECT 86.160000 95.575000 87.960000 96.825000 ;
        RECT 86.160000 87.435000 87.960000 88.685000 ;
        RECT 86.160000 79.295000 87.960000 80.545000 ;
        RECT 107.760000 95.575000 109.560000 96.825000 ;
        RECT 107.760000 87.435000 109.560000 88.685000 ;
        RECT 107.760000 79.295000 109.560000 80.545000 ;
        RECT 96.960000 111.855000 98.760000 113.105000 ;
        RECT 96.960000 103.715000 98.760000 104.965000 ;
        RECT 86.160000 111.855000 87.960000 113.105000 ;
        RECT 86.160000 103.715000 87.960000 104.965000 ;
        RECT 107.760000 111.855000 109.560000 113.105000 ;
        RECT 107.760000 103.715000 109.560000 104.965000 ;
        RECT 129.360000 87.435000 131.160000 88.685000 ;
        RECT 118.560000 87.435000 120.360000 88.685000 ;
        RECT 118.560000 79.295000 120.360000 80.545000 ;
        RECT 129.360000 79.295000 131.160000 80.545000 ;
        RECT 118.560000 95.575000 120.360000 96.825000 ;
        RECT 129.360000 95.575000 131.160000 96.825000 ;
        RECT 150.960000 95.575000 152.760000 96.825000 ;
        RECT 150.960000 87.435000 152.760000 88.685000 ;
        RECT 150.960000 79.295000 152.760000 80.545000 ;
        RECT 140.160000 95.575000 141.960000 96.825000 ;
        RECT 140.160000 87.435000 141.960000 88.685000 ;
        RECT 140.160000 79.295000 141.960000 80.545000 ;
        RECT 118.560000 103.715000 120.360000 104.965000 ;
        RECT 118.560000 111.855000 120.360000 113.105000 ;
        RECT 129.360000 103.715000 131.160000 104.965000 ;
        RECT 129.360000 111.855000 131.160000 113.105000 ;
        RECT 150.960000 111.855000 152.760000 113.105000 ;
        RECT 150.960000 103.715000 152.760000 104.965000 ;
        RECT 140.160000 111.855000 141.960000 113.105000 ;
        RECT 140.160000 103.715000 141.960000 104.965000 ;
        RECT 107.760000 136.275000 109.560000 137.525000 ;
        RECT 96.960000 136.275000 98.760000 137.525000 ;
        RECT 86.160000 136.275000 87.960000 137.525000 ;
        RECT 96.960000 128.135000 98.760000 129.385000 ;
        RECT 96.960000 119.995000 98.760000 121.245000 ;
        RECT 86.160000 128.135000 87.960000 129.385000 ;
        RECT 86.160000 119.995000 87.960000 121.245000 ;
        RECT 107.760000 128.135000 109.560000 129.385000 ;
        RECT 107.760000 119.995000 109.560000 121.245000 ;
        RECT 96.960000 152.555000 98.760000 153.805000 ;
        RECT 96.960000 144.415000 98.760000 145.665000 ;
        RECT 86.160000 152.555000 87.960000 153.805000 ;
        RECT 86.160000 144.415000 87.960000 145.665000 ;
        RECT 107.760000 152.555000 109.560000 153.805000 ;
        RECT 107.760000 144.415000 109.560000 145.665000 ;
        RECT 150.960000 136.275000 152.760000 137.525000 ;
        RECT 140.160000 136.275000 141.960000 137.525000 ;
        RECT 129.360000 136.275000 131.160000 137.525000 ;
        RECT 118.560000 136.275000 120.360000 137.525000 ;
        RECT 118.560000 119.995000 120.360000 121.245000 ;
        RECT 118.560000 128.135000 120.360000 129.385000 ;
        RECT 129.360000 119.995000 131.160000 121.245000 ;
        RECT 129.360000 128.135000 131.160000 129.385000 ;
        RECT 150.960000 128.135000 152.760000 129.385000 ;
        RECT 150.960000 119.995000 152.760000 121.245000 ;
        RECT 140.160000 128.135000 141.960000 129.385000 ;
        RECT 140.160000 119.995000 141.960000 121.245000 ;
        RECT 118.560000 144.415000 120.360000 145.665000 ;
        RECT 118.560000 152.555000 120.360000 153.805000 ;
        RECT 129.360000 144.415000 131.160000 145.665000 ;
        RECT 129.360000 152.555000 131.160000 153.805000 ;
        RECT 150.960000 152.555000 152.760000 153.805000 ;
        RECT 150.960000 144.415000 152.760000 145.665000 ;
        RECT 140.160000 152.555000 141.960000 153.805000 ;
        RECT 140.160000 144.415000 141.960000 145.665000 ;
        RECT 226.560000 38.595000 228.360000 39.845000 ;
        RECT 215.760000 38.595000 217.560000 39.845000 ;
        RECT 204.960000 38.595000 206.760000 39.845000 ;
        RECT 194.160000 38.595000 195.960000 39.845000 ;
        RECT 183.360000 38.595000 185.160000 39.845000 ;
        RECT 172.560000 38.595000 174.360000 39.845000 ;
        RECT 161.760000 38.595000 163.560000 39.845000 ;
        RECT 194.160000 30.455000 195.960000 31.705000 ;
        RECT 194.160000 22.315000 195.960000 23.565000 ;
        RECT 194.160000 14.175000 195.960000 15.425000 ;
        RECT 161.760000 14.175000 163.560000 15.425000 ;
        RECT 172.560000 14.175000 174.360000 15.425000 ;
        RECT 183.360000 14.175000 185.160000 15.425000 ;
        RECT 161.760000 22.315000 163.560000 23.565000 ;
        RECT 161.760000 30.455000 163.560000 31.705000 ;
        RECT 172.560000 22.315000 174.360000 23.565000 ;
        RECT 172.560000 30.455000 174.360000 31.705000 ;
        RECT 183.360000 22.315000 185.160000 23.565000 ;
        RECT 183.360000 30.455000 185.160000 31.705000 ;
        RECT 204.960000 14.175000 206.760000 15.425000 ;
        RECT 215.760000 14.175000 217.560000 15.425000 ;
        RECT 226.560000 14.175000 228.360000 15.425000 ;
        RECT 204.960000 22.315000 206.760000 23.565000 ;
        RECT 204.960000 30.455000 206.760000 31.705000 ;
        RECT 215.760000 22.315000 217.560000 23.565000 ;
        RECT 215.760000 30.455000 217.560000 31.705000 ;
        RECT 226.560000 22.315000 228.360000 23.565000 ;
        RECT 226.560000 30.455000 228.360000 31.705000 ;
        RECT 194.160000 71.155000 195.960000 72.405000 ;
        RECT 194.160000 63.015000 195.960000 64.265000 ;
        RECT 194.160000 54.875000 195.960000 56.125000 ;
        RECT 194.160000 46.735000 195.960000 47.985000 ;
        RECT 183.360000 54.875000 185.160000 56.125000 ;
        RECT 161.760000 46.735000 163.560000 47.985000 ;
        RECT 161.760000 54.875000 163.560000 56.125000 ;
        RECT 172.560000 46.735000 174.360000 47.985000 ;
        RECT 172.560000 54.875000 174.360000 56.125000 ;
        RECT 183.360000 46.735000 185.160000 47.985000 ;
        RECT 183.360000 71.155000 185.160000 72.405000 ;
        RECT 183.360000 63.015000 185.160000 64.265000 ;
        RECT 161.760000 63.015000 163.560000 64.265000 ;
        RECT 161.760000 71.155000 163.560000 72.405000 ;
        RECT 172.560000 63.015000 174.360000 64.265000 ;
        RECT 172.560000 71.155000 174.360000 72.405000 ;
        RECT 226.560000 54.875000 228.360000 56.125000 ;
        RECT 226.560000 46.735000 228.360000 47.985000 ;
        RECT 204.960000 46.735000 206.760000 47.985000 ;
        RECT 204.960000 54.875000 206.760000 56.125000 ;
        RECT 215.760000 46.735000 217.560000 47.985000 ;
        RECT 215.760000 54.875000 217.560000 56.125000 ;
        RECT 204.960000 71.155000 206.760000 72.405000 ;
        RECT 204.960000 63.015000 206.760000 64.265000 ;
        RECT 215.760000 63.015000 217.560000 64.265000 ;
        RECT 215.760000 71.155000 217.560000 72.405000 ;
        RECT 226.560000 63.015000 228.360000 64.265000 ;
        RECT 226.560000 71.155000 228.360000 72.405000 ;
        RECT 291.360000 38.595000 293.160000 39.845000 ;
        RECT 280.560000 38.595000 282.360000 39.845000 ;
        RECT 269.760000 38.595000 271.560000 39.845000 ;
        RECT 258.960000 38.595000 260.760000 39.845000 ;
        RECT 248.160000 38.595000 249.960000 39.845000 ;
        RECT 237.360000 38.595000 239.160000 39.845000 ;
        RECT 301.680000 38.595000 303.680000 39.845000 ;
        RECT 237.360000 14.175000 239.160000 15.425000 ;
        RECT 248.160000 14.175000 249.960000 15.425000 ;
        RECT 258.960000 14.175000 260.760000 15.425000 ;
        RECT 269.760000 14.175000 271.560000 15.425000 ;
        RECT 269.760000 30.455000 271.560000 31.705000 ;
        RECT 237.360000 22.315000 239.160000 23.565000 ;
        RECT 237.360000 30.455000 239.160000 31.705000 ;
        RECT 248.160000 22.315000 249.960000 23.565000 ;
        RECT 248.160000 30.455000 249.960000 31.705000 ;
        RECT 258.960000 22.315000 260.760000 23.565000 ;
        RECT 258.960000 30.455000 260.760000 31.705000 ;
        RECT 269.760000 22.315000 271.560000 23.565000 ;
        RECT 291.360000 14.175000 293.160000 15.425000 ;
        RECT 280.560000 14.175000 282.360000 15.425000 ;
        RECT 301.680000 14.175000 303.680000 15.425000 ;
        RECT 291.360000 30.455000 293.160000 31.705000 ;
        RECT 291.360000 22.315000 293.160000 23.565000 ;
        RECT 280.560000 30.455000 282.360000 31.705000 ;
        RECT 280.560000 22.315000 282.360000 23.565000 ;
        RECT 301.680000 30.455000 303.680000 31.705000 ;
        RECT 301.680000 22.315000 303.680000 23.565000 ;
        RECT 269.760000 54.875000 271.560000 56.125000 ;
        RECT 269.760000 46.735000 271.560000 47.985000 ;
        RECT 258.960000 54.875000 260.760000 56.125000 ;
        RECT 258.960000 46.735000 260.760000 47.985000 ;
        RECT 248.160000 54.875000 249.960000 56.125000 ;
        RECT 237.360000 46.735000 239.160000 47.985000 ;
        RECT 237.360000 54.875000 239.160000 56.125000 ;
        RECT 248.160000 46.735000 249.960000 47.985000 ;
        RECT 237.360000 71.155000 239.160000 72.405000 ;
        RECT 237.360000 63.015000 239.160000 64.265000 ;
        RECT 248.160000 63.015000 249.960000 64.265000 ;
        RECT 248.160000 71.155000 249.960000 72.405000 ;
        RECT 258.960000 63.015000 260.760000 64.265000 ;
        RECT 258.960000 71.155000 260.760000 72.405000 ;
        RECT 269.760000 63.015000 271.560000 64.265000 ;
        RECT 269.760000 71.155000 271.560000 72.405000 ;
        RECT 291.360000 54.875000 293.160000 56.125000 ;
        RECT 291.360000 46.735000 293.160000 47.985000 ;
        RECT 280.560000 54.875000 282.360000 56.125000 ;
        RECT 280.560000 46.735000 282.360000 47.985000 ;
        RECT 301.680000 46.735000 303.680000 47.985000 ;
        RECT 301.680000 54.875000 303.680000 56.125000 ;
        RECT 291.360000 71.155000 293.160000 72.405000 ;
        RECT 291.360000 63.015000 293.160000 64.265000 ;
        RECT 280.560000 63.015000 282.360000 64.265000 ;
        RECT 280.560000 71.155000 282.360000 72.405000 ;
        RECT 301.680000 63.015000 303.680000 64.265000 ;
        RECT 301.680000 71.155000 303.680000 72.405000 ;
        RECT 194.160000 111.855000 195.960000 113.105000 ;
        RECT 194.160000 103.715000 195.960000 104.965000 ;
        RECT 194.160000 95.575000 195.960000 96.825000 ;
        RECT 194.160000 87.435000 195.960000 88.685000 ;
        RECT 194.160000 79.295000 195.960000 80.545000 ;
        RECT 172.560000 95.575000 174.360000 96.825000 ;
        RECT 172.560000 87.435000 174.360000 88.685000 ;
        RECT 172.560000 79.295000 174.360000 80.545000 ;
        RECT 161.760000 79.295000 163.560000 80.545000 ;
        RECT 161.760000 87.435000 163.560000 88.685000 ;
        RECT 161.760000 95.575000 163.560000 96.825000 ;
        RECT 183.360000 95.575000 185.160000 96.825000 ;
        RECT 183.360000 87.435000 185.160000 88.685000 ;
        RECT 183.360000 79.295000 185.160000 80.545000 ;
        RECT 161.760000 103.715000 163.560000 104.965000 ;
        RECT 161.760000 111.855000 163.560000 113.105000 ;
        RECT 172.560000 103.715000 174.360000 104.965000 ;
        RECT 172.560000 111.855000 174.360000 113.105000 ;
        RECT 183.360000 103.715000 185.160000 104.965000 ;
        RECT 183.360000 111.855000 185.160000 113.105000 ;
        RECT 204.960000 95.575000 206.760000 96.825000 ;
        RECT 204.960000 87.435000 206.760000 88.685000 ;
        RECT 204.960000 79.295000 206.760000 80.545000 ;
        RECT 226.560000 87.435000 228.360000 88.685000 ;
        RECT 215.760000 87.435000 217.560000 88.685000 ;
        RECT 215.760000 79.295000 217.560000 80.545000 ;
        RECT 226.560000 79.295000 228.360000 80.545000 ;
        RECT 215.760000 95.575000 217.560000 96.825000 ;
        RECT 226.560000 95.575000 228.360000 96.825000 ;
        RECT 204.960000 111.855000 206.760000 113.105000 ;
        RECT 204.960000 103.715000 206.760000 104.965000 ;
        RECT 226.560000 111.855000 228.360000 113.105000 ;
        RECT 226.560000 103.715000 228.360000 104.965000 ;
        RECT 215.760000 111.855000 217.560000 113.105000 ;
        RECT 215.760000 103.715000 217.560000 104.965000 ;
        RECT 194.160000 152.555000 195.960000 153.805000 ;
        RECT 194.160000 144.415000 195.960000 145.665000 ;
        RECT 194.160000 136.275000 195.960000 137.525000 ;
        RECT 194.160000 128.135000 195.960000 129.385000 ;
        RECT 194.160000 119.995000 195.960000 121.245000 ;
        RECT 183.360000 136.275000 185.160000 137.525000 ;
        RECT 172.560000 136.275000 174.360000 137.525000 ;
        RECT 161.760000 136.275000 163.560000 137.525000 ;
        RECT 161.760000 119.995000 163.560000 121.245000 ;
        RECT 161.760000 128.135000 163.560000 129.385000 ;
        RECT 172.560000 119.995000 174.360000 121.245000 ;
        RECT 172.560000 128.135000 174.360000 129.385000 ;
        RECT 183.360000 119.995000 185.160000 121.245000 ;
        RECT 183.360000 128.135000 185.160000 129.385000 ;
        RECT 161.760000 144.415000 163.560000 145.665000 ;
        RECT 161.760000 152.555000 163.560000 153.805000 ;
        RECT 172.560000 144.415000 174.360000 145.665000 ;
        RECT 172.560000 152.555000 174.360000 153.805000 ;
        RECT 183.360000 144.415000 185.160000 145.665000 ;
        RECT 183.360000 152.555000 185.160000 153.805000 ;
        RECT 226.560000 136.275000 228.360000 137.525000 ;
        RECT 215.760000 136.275000 217.560000 137.525000 ;
        RECT 204.960000 136.275000 206.760000 137.525000 ;
        RECT 204.960000 128.135000 206.760000 129.385000 ;
        RECT 204.960000 119.995000 206.760000 121.245000 ;
        RECT 226.560000 128.135000 228.360000 129.385000 ;
        RECT 226.560000 119.995000 228.360000 121.245000 ;
        RECT 215.760000 128.135000 217.560000 129.385000 ;
        RECT 215.760000 119.995000 217.560000 121.245000 ;
        RECT 204.960000 152.555000 206.760000 153.805000 ;
        RECT 204.960000 144.415000 206.760000 145.665000 ;
        RECT 226.560000 152.555000 228.360000 153.805000 ;
        RECT 226.560000 144.415000 228.360000 145.665000 ;
        RECT 215.760000 152.555000 217.560000 153.805000 ;
        RECT 215.760000 144.415000 217.560000 145.665000 ;
        RECT 248.160000 95.575000 249.960000 96.825000 ;
        RECT 248.160000 87.435000 249.960000 88.685000 ;
        RECT 248.160000 79.295000 249.960000 80.545000 ;
        RECT 237.360000 95.575000 239.160000 96.825000 ;
        RECT 237.360000 87.435000 239.160000 88.685000 ;
        RECT 237.360000 79.295000 239.160000 80.545000 ;
        RECT 269.760000 95.575000 271.560000 96.825000 ;
        RECT 269.760000 87.435000 271.560000 88.685000 ;
        RECT 269.760000 79.295000 271.560000 80.545000 ;
        RECT 258.960000 95.575000 260.760000 96.825000 ;
        RECT 258.960000 87.435000 260.760000 88.685000 ;
        RECT 258.960000 79.295000 260.760000 80.545000 ;
        RECT 237.360000 103.715000 239.160000 104.965000 ;
        RECT 237.360000 111.855000 239.160000 113.105000 ;
        RECT 248.160000 103.715000 249.960000 104.965000 ;
        RECT 248.160000 111.855000 249.960000 113.105000 ;
        RECT 269.760000 111.855000 271.560000 113.105000 ;
        RECT 269.760000 103.715000 271.560000 104.965000 ;
        RECT 258.960000 111.855000 260.760000 113.105000 ;
        RECT 258.960000 103.715000 260.760000 104.965000 ;
        RECT 291.360000 95.575000 293.160000 96.825000 ;
        RECT 291.360000 87.435000 293.160000 88.685000 ;
        RECT 291.360000 79.295000 293.160000 80.545000 ;
        RECT 280.560000 95.575000 282.360000 96.825000 ;
        RECT 280.560000 87.435000 282.360000 88.685000 ;
        RECT 280.560000 79.295000 282.360000 80.545000 ;
        RECT 301.680000 79.295000 303.680000 80.545000 ;
        RECT 301.680000 87.435000 303.680000 88.685000 ;
        RECT 301.680000 95.575000 303.680000 96.825000 ;
        RECT 291.360000 111.855000 293.160000 113.105000 ;
        RECT 291.360000 103.715000 293.160000 104.965000 ;
        RECT 280.560000 111.855000 282.360000 113.105000 ;
        RECT 280.560000 103.715000 282.360000 104.965000 ;
        RECT 301.680000 103.715000 303.680000 104.965000 ;
        RECT 301.680000 111.855000 303.680000 113.105000 ;
        RECT 269.760000 136.275000 271.560000 137.525000 ;
        RECT 258.960000 136.275000 260.760000 137.525000 ;
        RECT 248.160000 136.275000 249.960000 137.525000 ;
        RECT 237.360000 136.275000 239.160000 137.525000 ;
        RECT 237.360000 119.995000 239.160000 121.245000 ;
        RECT 237.360000 128.135000 239.160000 129.385000 ;
        RECT 248.160000 119.995000 249.960000 121.245000 ;
        RECT 248.160000 128.135000 249.960000 129.385000 ;
        RECT 269.760000 128.135000 271.560000 129.385000 ;
        RECT 269.760000 119.995000 271.560000 121.245000 ;
        RECT 258.960000 128.135000 260.760000 129.385000 ;
        RECT 258.960000 119.995000 260.760000 121.245000 ;
        RECT 237.360000 144.415000 239.160000 145.665000 ;
        RECT 237.360000 152.555000 239.160000 153.805000 ;
        RECT 248.160000 144.415000 249.960000 145.665000 ;
        RECT 248.160000 152.555000 249.960000 153.805000 ;
        RECT 269.760000 152.555000 271.560000 153.805000 ;
        RECT 269.760000 144.415000 271.560000 145.665000 ;
        RECT 258.960000 152.555000 260.760000 153.805000 ;
        RECT 258.960000 144.415000 260.760000 145.665000 ;
        RECT 291.360000 136.275000 293.160000 137.525000 ;
        RECT 280.560000 136.275000 282.360000 137.525000 ;
        RECT 301.680000 136.275000 303.680000 137.525000 ;
        RECT 291.360000 128.135000 293.160000 129.385000 ;
        RECT 291.360000 119.995000 293.160000 121.245000 ;
        RECT 280.560000 128.135000 282.360000 129.385000 ;
        RECT 280.560000 119.995000 282.360000 121.245000 ;
        RECT 301.680000 119.995000 303.680000 121.245000 ;
        RECT 301.680000 128.135000 303.680000 129.385000 ;
        RECT 291.360000 152.555000 293.160000 153.805000 ;
        RECT 291.360000 144.415000 293.160000 145.665000 ;
        RECT 280.560000 152.555000 282.360000 153.805000 ;
        RECT 280.560000 144.415000 282.360000 145.665000 ;
        RECT 301.680000 144.415000 303.680000 145.665000 ;
        RECT 301.680000 152.555000 303.680000 153.805000 ;
        RECT 7.360000 160.695000 9.360000 161.945000 ;
        RECT 10.560000 160.695000 12.360000 161.945000 ;
        RECT 7.360000 168.835000 9.360000 170.085000 ;
        RECT 10.560000 168.835000 12.360000 170.085000 ;
        RECT 21.360000 160.695000 23.160000 161.945000 ;
        RECT 32.160000 160.695000 33.960000 161.945000 ;
        RECT 21.360000 168.835000 23.160000 170.085000 ;
        RECT 32.160000 168.835000 33.960000 170.085000 ;
        RECT 7.360000 176.975000 9.360000 178.225000 ;
        RECT 10.560000 176.975000 12.360000 178.225000 ;
        RECT 7.360000 193.255000 9.360000 194.505000 ;
        RECT 7.360000 185.115000 9.360000 186.365000 ;
        RECT 10.560000 185.115000 12.360000 186.365000 ;
        RECT 10.560000 193.255000 12.360000 194.505000 ;
        RECT 21.360000 176.975000 23.160000 178.225000 ;
        RECT 32.160000 176.975000 33.960000 178.225000 ;
        RECT 21.360000 185.115000 23.160000 186.365000 ;
        RECT 21.360000 193.255000 23.160000 194.505000 ;
        RECT 32.160000 185.115000 33.960000 186.365000 ;
        RECT 32.160000 193.255000 33.960000 194.505000 ;
        RECT 53.760000 168.835000 55.560000 170.085000 ;
        RECT 53.760000 160.695000 55.560000 161.945000 ;
        RECT 42.960000 168.835000 44.760000 170.085000 ;
        RECT 42.960000 160.695000 44.760000 161.945000 ;
        RECT 75.360000 168.835000 77.160000 170.085000 ;
        RECT 75.360000 160.695000 77.160000 161.945000 ;
        RECT 64.560000 168.835000 66.360000 170.085000 ;
        RECT 64.560000 160.695000 66.360000 161.945000 ;
        RECT 53.760000 193.255000 55.560000 194.505000 ;
        RECT 53.760000 185.115000 55.560000 186.365000 ;
        RECT 53.760000 176.975000 55.560000 178.225000 ;
        RECT 42.960000 193.255000 44.760000 194.505000 ;
        RECT 42.960000 185.115000 44.760000 186.365000 ;
        RECT 42.960000 176.975000 44.760000 178.225000 ;
        RECT 75.360000 193.255000 77.160000 194.505000 ;
        RECT 75.360000 185.115000 77.160000 186.365000 ;
        RECT 75.360000 176.975000 77.160000 178.225000 ;
        RECT 64.560000 193.255000 66.360000 194.505000 ;
        RECT 64.560000 185.115000 66.360000 186.365000 ;
        RECT 64.560000 176.975000 66.360000 178.225000 ;
        RECT 10.560000 209.535000 12.360000 210.785000 ;
        RECT 10.560000 201.395000 12.360000 202.645000 ;
        RECT 7.360000 201.395000 9.360000 202.645000 ;
        RECT 7.360000 209.535000 9.360000 210.785000 ;
        RECT 32.160000 209.535000 33.960000 210.785000 ;
        RECT 32.160000 201.395000 33.960000 202.645000 ;
        RECT 21.360000 209.535000 23.160000 210.785000 ;
        RECT 21.360000 201.395000 23.160000 202.645000 ;
        RECT 10.560000 225.815000 12.360000 227.065000 ;
        RECT 10.560000 217.675000 12.360000 218.925000 ;
        RECT 7.360000 217.675000 9.360000 218.925000 ;
        RECT 7.360000 225.815000 9.360000 227.065000 ;
        RECT 32.160000 225.815000 33.960000 227.065000 ;
        RECT 32.160000 217.675000 33.960000 218.925000 ;
        RECT 21.360000 225.815000 23.160000 227.065000 ;
        RECT 21.360000 217.675000 23.160000 218.925000 ;
        RECT 42.960000 201.395000 44.760000 202.645000 ;
        RECT 42.960000 209.535000 44.760000 210.785000 ;
        RECT 53.760000 201.395000 55.560000 202.645000 ;
        RECT 53.760000 209.535000 55.560000 210.785000 ;
        RECT 75.360000 209.535000 77.160000 210.785000 ;
        RECT 75.360000 201.395000 77.160000 202.645000 ;
        RECT 64.560000 209.535000 66.360000 210.785000 ;
        RECT 64.560000 201.395000 66.360000 202.645000 ;
        RECT 42.960000 217.675000 44.760000 218.925000 ;
        RECT 42.960000 225.815000 44.760000 227.065000 ;
        RECT 53.760000 217.675000 55.560000 218.925000 ;
        RECT 53.760000 225.815000 55.560000 227.065000 ;
        RECT 75.360000 225.815000 77.160000 227.065000 ;
        RECT 75.360000 217.675000 77.160000 218.925000 ;
        RECT 64.560000 225.815000 66.360000 227.065000 ;
        RECT 64.560000 217.675000 66.360000 218.925000 ;
        RECT 96.960000 168.835000 98.760000 170.085000 ;
        RECT 96.960000 160.695000 98.760000 161.945000 ;
        RECT 86.160000 168.835000 87.960000 170.085000 ;
        RECT 86.160000 160.695000 87.960000 161.945000 ;
        RECT 107.760000 168.835000 109.560000 170.085000 ;
        RECT 107.760000 160.695000 109.560000 161.945000 ;
        RECT 96.960000 193.255000 98.760000 194.505000 ;
        RECT 96.960000 185.115000 98.760000 186.365000 ;
        RECT 96.960000 176.975000 98.760000 178.225000 ;
        RECT 86.160000 193.255000 87.960000 194.505000 ;
        RECT 86.160000 185.115000 87.960000 186.365000 ;
        RECT 86.160000 176.975000 87.960000 178.225000 ;
        RECT 107.760000 193.255000 109.560000 194.505000 ;
        RECT 107.760000 185.115000 109.560000 186.365000 ;
        RECT 107.760000 176.975000 109.560000 178.225000 ;
        RECT 118.560000 160.695000 120.360000 161.945000 ;
        RECT 129.360000 160.695000 131.160000 161.945000 ;
        RECT 118.560000 168.835000 120.360000 170.085000 ;
        RECT 129.360000 168.835000 131.160000 170.085000 ;
        RECT 150.960000 168.835000 152.760000 170.085000 ;
        RECT 150.960000 160.695000 152.760000 161.945000 ;
        RECT 140.160000 168.835000 141.960000 170.085000 ;
        RECT 140.160000 160.695000 141.960000 161.945000 ;
        RECT 118.560000 176.975000 120.360000 178.225000 ;
        RECT 129.360000 176.975000 131.160000 178.225000 ;
        RECT 118.560000 185.115000 120.360000 186.365000 ;
        RECT 118.560000 193.255000 120.360000 194.505000 ;
        RECT 129.360000 185.115000 131.160000 186.365000 ;
        RECT 129.360000 193.255000 131.160000 194.505000 ;
        RECT 150.960000 193.255000 152.760000 194.505000 ;
        RECT 150.960000 185.115000 152.760000 186.365000 ;
        RECT 150.960000 176.975000 152.760000 178.225000 ;
        RECT 140.160000 193.255000 141.960000 194.505000 ;
        RECT 140.160000 185.115000 141.960000 186.365000 ;
        RECT 140.160000 176.975000 141.960000 178.225000 ;
        RECT 96.960000 209.535000 98.760000 210.785000 ;
        RECT 96.960000 201.395000 98.760000 202.645000 ;
        RECT 86.160000 209.535000 87.960000 210.785000 ;
        RECT 86.160000 201.395000 87.960000 202.645000 ;
        RECT 107.760000 209.535000 109.560000 210.785000 ;
        RECT 107.760000 201.395000 109.560000 202.645000 ;
        RECT 96.960000 225.815000 98.760000 227.065000 ;
        RECT 96.960000 217.675000 98.760000 218.925000 ;
        RECT 86.160000 225.815000 87.960000 227.065000 ;
        RECT 86.160000 217.675000 87.960000 218.925000 ;
        RECT 107.760000 225.815000 109.560000 227.065000 ;
        RECT 107.760000 217.675000 109.560000 218.925000 ;
        RECT 118.560000 201.395000 120.360000 202.645000 ;
        RECT 118.560000 209.535000 120.360000 210.785000 ;
        RECT 129.360000 201.395000 131.160000 202.645000 ;
        RECT 129.360000 209.535000 131.160000 210.785000 ;
        RECT 150.960000 209.535000 152.760000 210.785000 ;
        RECT 150.960000 201.395000 152.760000 202.645000 ;
        RECT 140.160000 209.535000 141.960000 210.785000 ;
        RECT 140.160000 201.395000 141.960000 202.645000 ;
        RECT 118.560000 217.675000 120.360000 218.925000 ;
        RECT 118.560000 225.815000 120.360000 227.065000 ;
        RECT 129.360000 217.675000 131.160000 218.925000 ;
        RECT 129.360000 225.815000 131.160000 227.065000 ;
        RECT 150.960000 225.815000 152.760000 227.065000 ;
        RECT 150.960000 217.675000 152.760000 218.925000 ;
        RECT 140.160000 225.815000 141.960000 227.065000 ;
        RECT 140.160000 217.675000 141.960000 218.925000 ;
        RECT 7.360000 242.095000 9.360000 243.345000 ;
        RECT 7.360000 233.955000 9.360000 235.205000 ;
        RECT 10.560000 233.955000 12.360000 235.205000 ;
        RECT 10.560000 242.095000 12.360000 243.345000 ;
        RECT 7.360000 250.235000 9.360000 251.485000 ;
        RECT 10.560000 250.235000 12.360000 251.485000 ;
        RECT 21.360000 233.955000 23.160000 235.205000 ;
        RECT 21.360000 242.095000 23.160000 243.345000 ;
        RECT 32.160000 233.955000 33.960000 235.205000 ;
        RECT 32.160000 242.095000 33.960000 243.345000 ;
        RECT 21.360000 250.235000 23.160000 251.485000 ;
        RECT 32.160000 250.235000 33.960000 251.485000 ;
        RECT 7.360000 258.375000 9.360000 259.625000 ;
        RECT 10.560000 258.375000 12.360000 259.625000 ;
        RECT 7.360000 266.515000 9.360000 267.765000 ;
        RECT 10.560000 266.515000 12.360000 267.765000 ;
        RECT 21.360000 258.375000 23.160000 259.625000 ;
        RECT 32.160000 258.375000 33.960000 259.625000 ;
        RECT 21.360000 266.515000 23.160000 267.765000 ;
        RECT 32.160000 266.515000 33.960000 267.765000 ;
        RECT 53.760000 250.235000 55.560000 251.485000 ;
        RECT 53.760000 242.095000 55.560000 243.345000 ;
        RECT 53.760000 233.955000 55.560000 235.205000 ;
        RECT 42.960000 250.235000 44.760000 251.485000 ;
        RECT 42.960000 242.095000 44.760000 243.345000 ;
        RECT 42.960000 233.955000 44.760000 235.205000 ;
        RECT 75.360000 250.235000 77.160000 251.485000 ;
        RECT 75.360000 242.095000 77.160000 243.345000 ;
        RECT 75.360000 233.955000 77.160000 235.205000 ;
        RECT 64.560000 250.235000 66.360000 251.485000 ;
        RECT 64.560000 242.095000 66.360000 243.345000 ;
        RECT 64.560000 233.955000 66.360000 235.205000 ;
        RECT 53.760000 266.515000 55.560000 267.765000 ;
        RECT 53.760000 258.375000 55.560000 259.625000 ;
        RECT 42.960000 266.515000 44.760000 267.765000 ;
        RECT 42.960000 258.375000 44.760000 259.625000 ;
        RECT 75.360000 266.515000 77.160000 267.765000 ;
        RECT 75.360000 258.375000 77.160000 259.625000 ;
        RECT 64.560000 266.515000 66.360000 267.765000 ;
        RECT 64.560000 258.375000 66.360000 259.625000 ;
        RECT 32.160000 290.935000 33.960000 292.185000 ;
        RECT 21.360000 290.935000 23.160000 292.185000 ;
        RECT 10.560000 290.935000 12.360000 292.185000 ;
        RECT 7.360000 290.935000 9.360000 292.185000 ;
        RECT 10.560000 282.795000 12.360000 284.045000 ;
        RECT 10.560000 274.655000 12.360000 275.905000 ;
        RECT 7.360000 274.655000 9.360000 275.905000 ;
        RECT 7.360000 282.795000 9.360000 284.045000 ;
        RECT 32.160000 282.795000 33.960000 284.045000 ;
        RECT 32.160000 274.655000 33.960000 275.905000 ;
        RECT 21.360000 282.795000 23.160000 284.045000 ;
        RECT 21.360000 274.655000 23.160000 275.905000 ;
        RECT 9.930000 299.075000 10.260000 299.445000 ;
        RECT 7.360000 299.535000 9.360000 299.865000 ;
        RECT 10.560000 299.075000 12.360000 299.865000 ;
        RECT 32.160000 299.075000 33.960000 299.865000 ;
        RECT 21.360000 299.075000 23.160000 299.865000 ;
        RECT 75.360000 290.935000 77.160000 292.185000 ;
        RECT 64.560000 290.935000 66.360000 292.185000 ;
        RECT 53.760000 290.935000 55.560000 292.185000 ;
        RECT 42.960000 290.935000 44.760000 292.185000 ;
        RECT 42.960000 274.655000 44.760000 275.905000 ;
        RECT 42.960000 282.795000 44.760000 284.045000 ;
        RECT 53.760000 274.655000 55.560000 275.905000 ;
        RECT 53.760000 282.795000 55.560000 284.045000 ;
        RECT 75.360000 282.795000 77.160000 284.045000 ;
        RECT 75.360000 274.655000 77.160000 275.905000 ;
        RECT 64.560000 282.795000 66.360000 284.045000 ;
        RECT 64.560000 274.655000 66.360000 275.905000 ;
        RECT 42.960000 299.075000 44.760000 299.865000 ;
        RECT 53.760000 299.075000 55.560000 299.865000 ;
        RECT 64.560000 299.075000 66.360000 299.865000 ;
        RECT 75.360000 299.075000 77.160000 299.865000 ;
        RECT 96.960000 250.235000 98.760000 251.485000 ;
        RECT 96.960000 242.095000 98.760000 243.345000 ;
        RECT 96.960000 233.955000 98.760000 235.205000 ;
        RECT 86.160000 250.235000 87.960000 251.485000 ;
        RECT 86.160000 242.095000 87.960000 243.345000 ;
        RECT 86.160000 233.955000 87.960000 235.205000 ;
        RECT 107.760000 250.235000 109.560000 251.485000 ;
        RECT 107.760000 242.095000 109.560000 243.345000 ;
        RECT 107.760000 233.955000 109.560000 235.205000 ;
        RECT 96.960000 266.515000 98.760000 267.765000 ;
        RECT 96.960000 258.375000 98.760000 259.625000 ;
        RECT 86.160000 266.515000 87.960000 267.765000 ;
        RECT 86.160000 258.375000 87.960000 259.625000 ;
        RECT 107.760000 266.515000 109.560000 267.765000 ;
        RECT 107.760000 258.375000 109.560000 259.625000 ;
        RECT 118.560000 233.955000 120.360000 235.205000 ;
        RECT 118.560000 242.095000 120.360000 243.345000 ;
        RECT 129.360000 233.955000 131.160000 235.205000 ;
        RECT 129.360000 242.095000 131.160000 243.345000 ;
        RECT 118.560000 250.235000 120.360000 251.485000 ;
        RECT 129.360000 250.235000 131.160000 251.485000 ;
        RECT 150.960000 250.235000 152.760000 251.485000 ;
        RECT 150.960000 242.095000 152.760000 243.345000 ;
        RECT 150.960000 233.955000 152.760000 235.205000 ;
        RECT 140.160000 250.235000 141.960000 251.485000 ;
        RECT 140.160000 242.095000 141.960000 243.345000 ;
        RECT 140.160000 233.955000 141.960000 235.205000 ;
        RECT 118.560000 258.375000 120.360000 259.625000 ;
        RECT 129.360000 258.375000 131.160000 259.625000 ;
        RECT 118.560000 266.515000 120.360000 267.765000 ;
        RECT 129.360000 266.515000 131.160000 267.765000 ;
        RECT 150.960000 266.515000 152.760000 267.765000 ;
        RECT 150.960000 258.375000 152.760000 259.625000 ;
        RECT 140.160000 266.515000 141.960000 267.765000 ;
        RECT 140.160000 258.375000 141.960000 259.625000 ;
        RECT 107.760000 290.935000 109.560000 292.185000 ;
        RECT 96.960000 290.935000 98.760000 292.185000 ;
        RECT 86.160000 290.935000 87.960000 292.185000 ;
        RECT 96.960000 282.795000 98.760000 284.045000 ;
        RECT 96.960000 274.655000 98.760000 275.905000 ;
        RECT 86.160000 282.795000 87.960000 284.045000 ;
        RECT 86.160000 274.655000 87.960000 275.905000 ;
        RECT 107.760000 282.795000 109.560000 284.045000 ;
        RECT 107.760000 274.655000 109.560000 275.905000 ;
        RECT 96.960000 299.075000 98.760000 299.865000 ;
        RECT 86.160000 299.075000 87.960000 299.865000 ;
        RECT 107.760000 299.075000 109.560000 299.865000 ;
        RECT 150.960000 290.935000 152.760000 292.185000 ;
        RECT 140.160000 290.935000 141.960000 292.185000 ;
        RECT 129.360000 290.935000 131.160000 292.185000 ;
        RECT 118.560000 290.935000 120.360000 292.185000 ;
        RECT 118.560000 274.655000 120.360000 275.905000 ;
        RECT 118.560000 282.795000 120.360000 284.045000 ;
        RECT 129.360000 274.655000 131.160000 275.905000 ;
        RECT 129.360000 282.795000 131.160000 284.045000 ;
        RECT 150.960000 282.795000 152.760000 284.045000 ;
        RECT 150.960000 274.655000 152.760000 275.905000 ;
        RECT 140.160000 282.795000 141.960000 284.045000 ;
        RECT 140.160000 274.655000 141.960000 275.905000 ;
        RECT 118.560000 299.075000 120.360000 299.865000 ;
        RECT 129.360000 299.075000 131.160000 299.865000 ;
        RECT 140.160000 299.075000 141.960000 299.865000 ;
        RECT 150.960000 299.075000 152.760000 299.865000 ;
        RECT 194.160000 193.255000 195.960000 194.505000 ;
        RECT 194.160000 185.115000 195.960000 186.365000 ;
        RECT 194.160000 176.975000 195.960000 178.225000 ;
        RECT 194.160000 168.835000 195.960000 170.085000 ;
        RECT 194.160000 160.695000 195.960000 161.945000 ;
        RECT 172.560000 168.835000 174.360000 170.085000 ;
        RECT 172.560000 160.695000 174.360000 161.945000 ;
        RECT 161.760000 168.835000 163.560000 170.085000 ;
        RECT 161.760000 160.695000 163.560000 161.945000 ;
        RECT 183.360000 168.835000 185.160000 170.085000 ;
        RECT 183.360000 160.695000 185.160000 161.945000 ;
        RECT 172.560000 193.255000 174.360000 194.505000 ;
        RECT 172.560000 185.115000 174.360000 186.365000 ;
        RECT 172.560000 176.975000 174.360000 178.225000 ;
        RECT 161.760000 176.975000 163.560000 178.225000 ;
        RECT 161.760000 185.115000 163.560000 186.365000 ;
        RECT 161.760000 193.255000 163.560000 194.505000 ;
        RECT 183.360000 193.255000 185.160000 194.505000 ;
        RECT 183.360000 185.115000 185.160000 186.365000 ;
        RECT 183.360000 176.975000 185.160000 178.225000 ;
        RECT 204.960000 168.835000 206.760000 170.085000 ;
        RECT 204.960000 160.695000 206.760000 161.945000 ;
        RECT 215.760000 160.695000 217.560000 161.945000 ;
        RECT 226.560000 160.695000 228.360000 161.945000 ;
        RECT 215.760000 168.835000 217.560000 170.085000 ;
        RECT 226.560000 168.835000 228.360000 170.085000 ;
        RECT 204.960000 193.255000 206.760000 194.505000 ;
        RECT 204.960000 185.115000 206.760000 186.365000 ;
        RECT 204.960000 176.975000 206.760000 178.225000 ;
        RECT 215.760000 176.975000 217.560000 178.225000 ;
        RECT 226.560000 176.975000 228.360000 178.225000 ;
        RECT 215.760000 185.115000 217.560000 186.365000 ;
        RECT 215.760000 193.255000 217.560000 194.505000 ;
        RECT 226.560000 185.115000 228.360000 186.365000 ;
        RECT 226.560000 193.255000 228.360000 194.505000 ;
        RECT 194.160000 225.815000 195.960000 227.065000 ;
        RECT 194.160000 217.675000 195.960000 218.925000 ;
        RECT 194.160000 209.535000 195.960000 210.785000 ;
        RECT 194.160000 201.395000 195.960000 202.645000 ;
        RECT 161.760000 201.395000 163.560000 202.645000 ;
        RECT 161.760000 209.535000 163.560000 210.785000 ;
        RECT 172.560000 201.395000 174.360000 202.645000 ;
        RECT 172.560000 209.535000 174.360000 210.785000 ;
        RECT 183.360000 201.395000 185.160000 202.645000 ;
        RECT 183.360000 209.535000 185.160000 210.785000 ;
        RECT 161.760000 217.675000 163.560000 218.925000 ;
        RECT 161.760000 225.815000 163.560000 227.065000 ;
        RECT 172.560000 217.675000 174.360000 218.925000 ;
        RECT 172.560000 225.815000 174.360000 227.065000 ;
        RECT 183.360000 217.675000 185.160000 218.925000 ;
        RECT 183.360000 225.815000 185.160000 227.065000 ;
        RECT 204.960000 209.535000 206.760000 210.785000 ;
        RECT 204.960000 201.395000 206.760000 202.645000 ;
        RECT 226.560000 209.535000 228.360000 210.785000 ;
        RECT 226.560000 201.395000 228.360000 202.645000 ;
        RECT 215.760000 209.535000 217.560000 210.785000 ;
        RECT 215.760000 201.395000 217.560000 202.645000 ;
        RECT 204.960000 225.815000 206.760000 227.065000 ;
        RECT 204.960000 217.675000 206.760000 218.925000 ;
        RECT 226.560000 225.815000 228.360000 227.065000 ;
        RECT 226.560000 217.675000 228.360000 218.925000 ;
        RECT 215.760000 225.815000 217.560000 227.065000 ;
        RECT 215.760000 217.675000 217.560000 218.925000 ;
        RECT 248.160000 168.835000 249.960000 170.085000 ;
        RECT 248.160000 160.695000 249.960000 161.945000 ;
        RECT 237.360000 168.835000 239.160000 170.085000 ;
        RECT 237.360000 160.695000 239.160000 161.945000 ;
        RECT 269.760000 168.835000 271.560000 170.085000 ;
        RECT 269.760000 160.695000 271.560000 161.945000 ;
        RECT 258.960000 168.835000 260.760000 170.085000 ;
        RECT 258.960000 160.695000 260.760000 161.945000 ;
        RECT 248.160000 193.255000 249.960000 194.505000 ;
        RECT 248.160000 185.115000 249.960000 186.365000 ;
        RECT 248.160000 176.975000 249.960000 178.225000 ;
        RECT 237.360000 193.255000 239.160000 194.505000 ;
        RECT 237.360000 185.115000 239.160000 186.365000 ;
        RECT 237.360000 176.975000 239.160000 178.225000 ;
        RECT 269.760000 193.255000 271.560000 194.505000 ;
        RECT 269.760000 185.115000 271.560000 186.365000 ;
        RECT 269.760000 176.975000 271.560000 178.225000 ;
        RECT 258.960000 193.255000 260.760000 194.505000 ;
        RECT 258.960000 185.115000 260.760000 186.365000 ;
        RECT 258.960000 176.975000 260.760000 178.225000 ;
        RECT 291.360000 168.835000 293.160000 170.085000 ;
        RECT 291.360000 160.695000 293.160000 161.945000 ;
        RECT 280.560000 168.835000 282.360000 170.085000 ;
        RECT 280.560000 160.695000 282.360000 161.945000 ;
        RECT 301.680000 168.835000 303.680000 170.085000 ;
        RECT 301.680000 160.695000 303.680000 161.945000 ;
        RECT 291.360000 193.255000 293.160000 194.505000 ;
        RECT 291.360000 185.115000 293.160000 186.365000 ;
        RECT 291.360000 176.975000 293.160000 178.225000 ;
        RECT 280.560000 193.255000 282.360000 194.505000 ;
        RECT 280.560000 185.115000 282.360000 186.365000 ;
        RECT 280.560000 176.975000 282.360000 178.225000 ;
        RECT 301.680000 176.975000 303.680000 178.225000 ;
        RECT 301.680000 185.115000 303.680000 186.365000 ;
        RECT 301.680000 193.255000 303.680000 194.505000 ;
        RECT 237.360000 201.395000 239.160000 202.645000 ;
        RECT 237.360000 209.535000 239.160000 210.785000 ;
        RECT 248.160000 201.395000 249.960000 202.645000 ;
        RECT 248.160000 209.535000 249.960000 210.785000 ;
        RECT 269.760000 209.535000 271.560000 210.785000 ;
        RECT 269.760000 201.395000 271.560000 202.645000 ;
        RECT 258.960000 209.535000 260.760000 210.785000 ;
        RECT 258.960000 201.395000 260.760000 202.645000 ;
        RECT 237.360000 217.675000 239.160000 218.925000 ;
        RECT 237.360000 225.815000 239.160000 227.065000 ;
        RECT 248.160000 217.675000 249.960000 218.925000 ;
        RECT 248.160000 225.815000 249.960000 227.065000 ;
        RECT 269.760000 225.815000 271.560000 227.065000 ;
        RECT 269.760000 217.675000 271.560000 218.925000 ;
        RECT 258.960000 225.815000 260.760000 227.065000 ;
        RECT 258.960000 217.675000 260.760000 218.925000 ;
        RECT 291.360000 209.535000 293.160000 210.785000 ;
        RECT 291.360000 201.395000 293.160000 202.645000 ;
        RECT 280.560000 209.535000 282.360000 210.785000 ;
        RECT 280.560000 201.395000 282.360000 202.645000 ;
        RECT 301.680000 201.395000 303.680000 202.645000 ;
        RECT 301.680000 209.535000 303.680000 210.785000 ;
        RECT 291.360000 225.815000 293.160000 227.065000 ;
        RECT 291.360000 217.675000 293.160000 218.925000 ;
        RECT 280.560000 225.815000 282.360000 227.065000 ;
        RECT 280.560000 217.675000 282.360000 218.925000 ;
        RECT 301.680000 217.675000 303.680000 218.925000 ;
        RECT 301.680000 225.815000 303.680000 227.065000 ;
        RECT 194.160000 266.515000 195.960000 267.765000 ;
        RECT 194.160000 258.375000 195.960000 259.625000 ;
        RECT 194.160000 250.235000 195.960000 251.485000 ;
        RECT 194.160000 242.095000 195.960000 243.345000 ;
        RECT 194.160000 233.955000 195.960000 235.205000 ;
        RECT 172.560000 250.235000 174.360000 251.485000 ;
        RECT 172.560000 242.095000 174.360000 243.345000 ;
        RECT 172.560000 233.955000 174.360000 235.205000 ;
        RECT 161.760000 233.955000 163.560000 235.205000 ;
        RECT 161.760000 242.095000 163.560000 243.345000 ;
        RECT 161.760000 250.235000 163.560000 251.485000 ;
        RECT 183.360000 250.235000 185.160000 251.485000 ;
        RECT 183.360000 242.095000 185.160000 243.345000 ;
        RECT 183.360000 233.955000 185.160000 235.205000 ;
        RECT 172.560000 266.515000 174.360000 267.765000 ;
        RECT 172.560000 258.375000 174.360000 259.625000 ;
        RECT 161.760000 266.515000 163.560000 267.765000 ;
        RECT 161.760000 258.375000 163.560000 259.625000 ;
        RECT 183.360000 266.515000 185.160000 267.765000 ;
        RECT 183.360000 258.375000 185.160000 259.625000 ;
        RECT 204.960000 250.235000 206.760000 251.485000 ;
        RECT 204.960000 242.095000 206.760000 243.345000 ;
        RECT 204.960000 233.955000 206.760000 235.205000 ;
        RECT 215.760000 233.955000 217.560000 235.205000 ;
        RECT 215.760000 242.095000 217.560000 243.345000 ;
        RECT 226.560000 233.955000 228.360000 235.205000 ;
        RECT 226.560000 242.095000 228.360000 243.345000 ;
        RECT 215.760000 250.235000 217.560000 251.485000 ;
        RECT 226.560000 250.235000 228.360000 251.485000 ;
        RECT 204.960000 266.515000 206.760000 267.765000 ;
        RECT 204.960000 258.375000 206.760000 259.625000 ;
        RECT 215.760000 258.375000 217.560000 259.625000 ;
        RECT 226.560000 258.375000 228.360000 259.625000 ;
        RECT 215.760000 266.515000 217.560000 267.765000 ;
        RECT 226.560000 266.515000 228.360000 267.765000 ;
        RECT 194.160000 299.075000 195.960000 299.865000 ;
        RECT 194.160000 290.935000 195.960000 292.185000 ;
        RECT 194.160000 282.795000 195.960000 284.045000 ;
        RECT 194.160000 274.655000 195.960000 275.905000 ;
        RECT 183.360000 290.935000 185.160000 292.185000 ;
        RECT 172.560000 290.935000 174.360000 292.185000 ;
        RECT 161.760000 290.935000 163.560000 292.185000 ;
        RECT 161.760000 274.655000 163.560000 275.905000 ;
        RECT 161.760000 282.795000 163.560000 284.045000 ;
        RECT 172.560000 274.655000 174.360000 275.905000 ;
        RECT 172.560000 282.795000 174.360000 284.045000 ;
        RECT 183.360000 274.655000 185.160000 275.905000 ;
        RECT 183.360000 282.795000 185.160000 284.045000 ;
        RECT 183.360000 299.075000 185.160000 299.865000 ;
        RECT 172.560000 299.075000 174.360000 299.865000 ;
        RECT 161.760000 299.075000 163.560000 299.865000 ;
        RECT 226.560000 290.935000 228.360000 292.185000 ;
        RECT 215.760000 290.935000 217.560000 292.185000 ;
        RECT 204.960000 290.935000 206.760000 292.185000 ;
        RECT 204.960000 282.795000 206.760000 284.045000 ;
        RECT 204.960000 274.655000 206.760000 275.905000 ;
        RECT 226.560000 282.795000 228.360000 284.045000 ;
        RECT 226.560000 274.655000 228.360000 275.905000 ;
        RECT 215.760000 282.795000 217.560000 284.045000 ;
        RECT 215.760000 274.655000 217.560000 275.905000 ;
        RECT 204.960000 299.075000 206.760000 299.865000 ;
        RECT 215.760000 299.075000 217.560000 299.865000 ;
        RECT 226.560000 299.075000 228.360000 299.865000 ;
        RECT 248.160000 250.235000 249.960000 251.485000 ;
        RECT 248.160000 242.095000 249.960000 243.345000 ;
        RECT 248.160000 233.955000 249.960000 235.205000 ;
        RECT 237.360000 250.235000 239.160000 251.485000 ;
        RECT 237.360000 242.095000 239.160000 243.345000 ;
        RECT 237.360000 233.955000 239.160000 235.205000 ;
        RECT 269.760000 250.235000 271.560000 251.485000 ;
        RECT 269.760000 242.095000 271.560000 243.345000 ;
        RECT 269.760000 233.955000 271.560000 235.205000 ;
        RECT 258.960000 250.235000 260.760000 251.485000 ;
        RECT 258.960000 242.095000 260.760000 243.345000 ;
        RECT 258.960000 233.955000 260.760000 235.205000 ;
        RECT 248.160000 266.515000 249.960000 267.765000 ;
        RECT 248.160000 258.375000 249.960000 259.625000 ;
        RECT 237.360000 266.515000 239.160000 267.765000 ;
        RECT 237.360000 258.375000 239.160000 259.625000 ;
        RECT 269.760000 266.515000 271.560000 267.765000 ;
        RECT 269.760000 258.375000 271.560000 259.625000 ;
        RECT 258.960000 266.515000 260.760000 267.765000 ;
        RECT 258.960000 258.375000 260.760000 259.625000 ;
        RECT 291.360000 250.235000 293.160000 251.485000 ;
        RECT 291.360000 242.095000 293.160000 243.345000 ;
        RECT 291.360000 233.955000 293.160000 235.205000 ;
        RECT 280.560000 250.235000 282.360000 251.485000 ;
        RECT 280.560000 242.095000 282.360000 243.345000 ;
        RECT 280.560000 233.955000 282.360000 235.205000 ;
        RECT 301.680000 233.955000 303.680000 235.205000 ;
        RECT 301.680000 242.095000 303.680000 243.345000 ;
        RECT 301.680000 250.235000 303.680000 251.485000 ;
        RECT 291.360000 266.515000 293.160000 267.765000 ;
        RECT 291.360000 258.375000 293.160000 259.625000 ;
        RECT 280.560000 266.515000 282.360000 267.765000 ;
        RECT 280.560000 258.375000 282.360000 259.625000 ;
        RECT 301.680000 266.515000 303.680000 267.765000 ;
        RECT 301.680000 258.375000 303.680000 259.625000 ;
        RECT 269.760000 290.935000 271.560000 292.185000 ;
        RECT 258.960000 290.935000 260.760000 292.185000 ;
        RECT 248.160000 290.935000 249.960000 292.185000 ;
        RECT 237.360000 290.935000 239.160000 292.185000 ;
        RECT 237.360000 274.655000 239.160000 275.905000 ;
        RECT 237.360000 282.795000 239.160000 284.045000 ;
        RECT 248.160000 274.655000 249.960000 275.905000 ;
        RECT 248.160000 282.795000 249.960000 284.045000 ;
        RECT 269.760000 282.795000 271.560000 284.045000 ;
        RECT 269.760000 274.655000 271.560000 275.905000 ;
        RECT 258.960000 282.795000 260.760000 284.045000 ;
        RECT 258.960000 274.655000 260.760000 275.905000 ;
        RECT 237.360000 299.075000 239.160000 299.865000 ;
        RECT 248.160000 299.075000 249.960000 299.865000 ;
        RECT 258.960000 299.075000 260.760000 299.865000 ;
        RECT 269.760000 299.075000 271.560000 299.865000 ;
        RECT 291.360000 290.935000 293.160000 292.185000 ;
        RECT 280.560000 290.935000 282.360000 292.185000 ;
        RECT 301.680000 290.935000 303.680000 292.185000 ;
        RECT 291.360000 282.795000 293.160000 284.045000 ;
        RECT 291.360000 274.655000 293.160000 275.905000 ;
        RECT 280.560000 282.795000 282.360000 284.045000 ;
        RECT 280.560000 274.655000 282.360000 275.905000 ;
        RECT 301.680000 274.655000 303.680000 275.905000 ;
        RECT 301.680000 282.795000 303.680000 284.045000 ;
        RECT 291.360000 299.075000 293.160000 299.865000 ;
        RECT 280.560000 299.075000 282.360000 299.865000 ;
        RECT 300.780000 298.895000 301.110000 299.625000 ;
        RECT 301.680000 299.535000 303.680000 299.865000 ;
      LAYER met3 ;
        RECT 0.000000 7.530000 311.040000 9.530000 ;
        RECT 0.000000 300.900000 311.040000 302.900000 ;
        RECT 9.975000 299.075000 10.095000 299.445000 ;
        RECT 300.945000 299.075000 301.055000 299.445000 ;
        RECT 9.930000 299.075000 10.260000 299.445000 ;
        RECT 300.780000 298.895000 301.110000 299.625000 ;
        RECT 7.360000 38.595000 9.360000 39.845000 ;
        RECT 10.560000 38.595000 12.360000 39.845000 ;
        RECT 21.360000 38.595000 23.160000 39.845000 ;
        RECT 32.160000 38.595000 33.960000 39.845000 ;
        RECT 42.960000 38.595000 44.760000 39.845000 ;
        RECT 53.760000 38.595000 55.560000 39.845000 ;
        RECT 64.560000 38.595000 66.360000 39.845000 ;
        RECT 75.360000 38.595000 77.160000 39.845000 ;
        RECT 32.160000 14.175000 33.960000 15.425000 ;
        RECT 21.360000 14.175000 23.160000 15.425000 ;
        RECT 10.560000 14.175000 12.360000 15.425000 ;
        RECT 7.360000 14.175000 9.360000 15.425000 ;
        RECT 7.360000 22.315000 9.360000 23.565000 ;
        RECT 7.360000 30.455000 9.360000 31.705000 ;
        RECT 10.560000 22.315000 12.360000 23.565000 ;
        RECT 10.560000 30.455000 12.360000 31.705000 ;
        RECT 21.360000 22.315000 23.160000 23.565000 ;
        RECT 21.360000 30.455000 23.160000 31.705000 ;
        RECT 32.160000 22.315000 33.960000 23.565000 ;
        RECT 32.160000 30.455000 33.960000 31.705000 ;
        RECT 42.960000 14.175000 44.760000 15.425000 ;
        RECT 53.760000 14.175000 55.560000 15.425000 ;
        RECT 64.560000 14.175000 66.360000 15.425000 ;
        RECT 75.360000 14.175000 77.160000 15.425000 ;
        RECT 42.960000 22.315000 44.760000 23.565000 ;
        RECT 42.960000 30.455000 44.760000 31.705000 ;
        RECT 53.760000 22.315000 55.560000 23.565000 ;
        RECT 53.760000 30.455000 55.560000 31.705000 ;
        RECT 64.560000 22.315000 66.360000 23.565000 ;
        RECT 64.560000 30.455000 66.360000 31.705000 ;
        RECT 75.360000 22.315000 77.160000 23.565000 ;
        RECT 75.360000 30.455000 77.160000 31.705000 ;
        RECT 7.360000 46.735000 9.360000 47.985000 ;
        RECT 7.360000 54.875000 9.360000 56.125000 ;
        RECT 10.560000 46.735000 12.360000 47.985000 ;
        RECT 10.560000 54.875000 12.360000 56.125000 ;
        RECT 21.360000 46.735000 23.160000 47.985000 ;
        RECT 21.360000 54.875000 23.160000 56.125000 ;
        RECT 32.160000 46.735000 33.960000 47.985000 ;
        RECT 32.160000 54.875000 33.960000 56.125000 ;
        RECT 7.360000 63.015000 9.360000 64.265000 ;
        RECT 7.360000 71.155000 9.360000 72.405000 ;
        RECT 10.560000 63.015000 12.360000 64.265000 ;
        RECT 10.560000 71.155000 12.360000 72.405000 ;
        RECT 21.360000 63.015000 23.160000 64.265000 ;
        RECT 21.360000 71.155000 23.160000 72.405000 ;
        RECT 32.160000 63.015000 33.960000 64.265000 ;
        RECT 32.160000 71.155000 33.960000 72.405000 ;
        RECT 42.960000 46.735000 44.760000 47.985000 ;
        RECT 42.960000 54.875000 44.760000 56.125000 ;
        RECT 53.760000 46.735000 55.560000 47.985000 ;
        RECT 53.760000 54.875000 55.560000 56.125000 ;
        RECT 64.560000 46.735000 66.360000 47.985000 ;
        RECT 64.560000 54.875000 66.360000 56.125000 ;
        RECT 75.360000 46.735000 77.160000 47.985000 ;
        RECT 75.360000 54.875000 77.160000 56.125000 ;
        RECT 53.760000 71.155000 55.560000 72.405000 ;
        RECT 53.760000 63.015000 55.560000 64.265000 ;
        RECT 42.960000 71.155000 44.760000 72.405000 ;
        RECT 42.960000 63.015000 44.760000 64.265000 ;
        RECT 75.360000 71.155000 77.160000 72.405000 ;
        RECT 75.360000 63.015000 77.160000 64.265000 ;
        RECT 64.560000 71.155000 66.360000 72.405000 ;
        RECT 64.560000 63.015000 66.360000 64.265000 ;
        RECT 150.960000 38.595000 152.760000 39.845000 ;
        RECT 140.160000 38.595000 141.960000 39.845000 ;
        RECT 129.360000 38.595000 131.160000 39.845000 ;
        RECT 118.560000 38.595000 120.360000 39.845000 ;
        RECT 107.760000 38.595000 109.560000 39.845000 ;
        RECT 96.960000 38.595000 98.760000 39.845000 ;
        RECT 86.160000 38.595000 87.960000 39.845000 ;
        RECT 107.760000 14.175000 109.560000 15.425000 ;
        RECT 96.960000 14.175000 98.760000 15.425000 ;
        RECT 86.160000 14.175000 87.960000 15.425000 ;
        RECT 107.760000 30.455000 109.560000 31.705000 ;
        RECT 107.760000 22.315000 109.560000 23.565000 ;
        RECT 96.960000 30.455000 98.760000 31.705000 ;
        RECT 96.960000 22.315000 98.760000 23.565000 ;
        RECT 86.160000 30.455000 87.960000 31.705000 ;
        RECT 86.160000 22.315000 87.960000 23.565000 ;
        RECT 140.160000 14.175000 141.960000 15.425000 ;
        RECT 129.360000 14.175000 131.160000 15.425000 ;
        RECT 118.560000 14.175000 120.360000 15.425000 ;
        RECT 150.960000 14.175000 152.760000 15.425000 ;
        RECT 129.360000 30.455000 131.160000 31.705000 ;
        RECT 129.360000 22.315000 131.160000 23.565000 ;
        RECT 118.560000 30.455000 120.360000 31.705000 ;
        RECT 118.560000 22.315000 120.360000 23.565000 ;
        RECT 140.160000 22.315000 141.960000 23.565000 ;
        RECT 140.160000 30.455000 141.960000 31.705000 ;
        RECT 150.960000 22.315000 152.760000 23.565000 ;
        RECT 150.960000 30.455000 152.760000 31.705000 ;
        RECT 107.760000 46.735000 109.560000 47.985000 ;
        RECT 96.960000 54.875000 98.760000 56.125000 ;
        RECT 96.960000 46.735000 98.760000 47.985000 ;
        RECT 86.160000 54.875000 87.960000 56.125000 ;
        RECT 86.160000 46.735000 87.960000 47.985000 ;
        RECT 107.760000 54.875000 109.560000 56.125000 ;
        RECT 96.960000 71.155000 98.760000 72.405000 ;
        RECT 96.960000 63.015000 98.760000 64.265000 ;
        RECT 86.160000 63.015000 87.960000 64.265000 ;
        RECT 86.160000 71.155000 87.960000 72.405000 ;
        RECT 107.760000 71.155000 109.560000 72.405000 ;
        RECT 107.760000 63.015000 109.560000 64.265000 ;
        RECT 118.560000 46.735000 120.360000 47.985000 ;
        RECT 118.560000 54.875000 120.360000 56.125000 ;
        RECT 129.360000 46.735000 131.160000 47.985000 ;
        RECT 129.360000 54.875000 131.160000 56.125000 ;
        RECT 140.160000 46.735000 141.960000 47.985000 ;
        RECT 140.160000 54.875000 141.960000 56.125000 ;
        RECT 150.960000 46.735000 152.760000 47.985000 ;
        RECT 150.960000 54.875000 152.760000 56.125000 ;
        RECT 129.360000 71.155000 131.160000 72.405000 ;
        RECT 129.360000 63.015000 131.160000 64.265000 ;
        RECT 118.560000 71.155000 120.360000 72.405000 ;
        RECT 118.560000 63.015000 120.360000 64.265000 ;
        RECT 150.960000 71.155000 152.760000 72.405000 ;
        RECT 150.960000 63.015000 152.760000 64.265000 ;
        RECT 140.160000 71.155000 141.960000 72.405000 ;
        RECT 140.160000 63.015000 141.960000 64.265000 ;
        RECT 10.560000 87.435000 12.360000 88.685000 ;
        RECT 7.360000 87.435000 9.360000 88.685000 ;
        RECT 7.360000 79.295000 9.360000 80.545000 ;
        RECT 10.560000 79.295000 12.360000 80.545000 ;
        RECT 7.360000 95.575000 9.360000 96.825000 ;
        RECT 10.560000 95.575000 12.360000 96.825000 ;
        RECT 32.160000 87.435000 33.960000 88.685000 ;
        RECT 21.360000 87.435000 23.160000 88.685000 ;
        RECT 21.360000 79.295000 23.160000 80.545000 ;
        RECT 32.160000 79.295000 33.960000 80.545000 ;
        RECT 21.360000 95.575000 23.160000 96.825000 ;
        RECT 32.160000 95.575000 33.960000 96.825000 ;
        RECT 10.560000 111.855000 12.360000 113.105000 ;
        RECT 10.560000 103.715000 12.360000 104.965000 ;
        RECT 7.360000 103.715000 9.360000 104.965000 ;
        RECT 7.360000 111.855000 9.360000 113.105000 ;
        RECT 32.160000 111.855000 33.960000 113.105000 ;
        RECT 32.160000 103.715000 33.960000 104.965000 ;
        RECT 21.360000 111.855000 23.160000 113.105000 ;
        RECT 21.360000 103.715000 23.160000 104.965000 ;
        RECT 42.960000 79.295000 44.760000 80.545000 ;
        RECT 42.960000 87.435000 44.760000 88.685000 ;
        RECT 42.960000 95.575000 44.760000 96.825000 ;
        RECT 53.760000 79.295000 55.560000 80.545000 ;
        RECT 53.760000 87.435000 55.560000 88.685000 ;
        RECT 53.760000 95.575000 55.560000 96.825000 ;
        RECT 64.560000 79.295000 66.360000 80.545000 ;
        RECT 64.560000 87.435000 66.360000 88.685000 ;
        RECT 64.560000 95.575000 66.360000 96.825000 ;
        RECT 75.360000 79.295000 77.160000 80.545000 ;
        RECT 75.360000 87.435000 77.160000 88.685000 ;
        RECT 75.360000 95.575000 77.160000 96.825000 ;
        RECT 42.960000 103.715000 44.760000 104.965000 ;
        RECT 42.960000 111.855000 44.760000 113.105000 ;
        RECT 53.760000 103.715000 55.560000 104.965000 ;
        RECT 53.760000 111.855000 55.560000 113.105000 ;
        RECT 64.560000 103.715000 66.360000 104.965000 ;
        RECT 64.560000 111.855000 66.360000 113.105000 ;
        RECT 75.360000 103.715000 77.160000 104.965000 ;
        RECT 75.360000 111.855000 77.160000 113.105000 ;
        RECT 32.160000 136.275000 33.960000 137.525000 ;
        RECT 21.360000 136.275000 23.160000 137.525000 ;
        RECT 10.560000 136.275000 12.360000 137.525000 ;
        RECT 7.360000 136.275000 9.360000 137.525000 ;
        RECT 10.560000 128.135000 12.360000 129.385000 ;
        RECT 10.560000 119.995000 12.360000 121.245000 ;
        RECT 7.360000 119.995000 9.360000 121.245000 ;
        RECT 7.360000 128.135000 9.360000 129.385000 ;
        RECT 32.160000 128.135000 33.960000 129.385000 ;
        RECT 32.160000 119.995000 33.960000 121.245000 ;
        RECT 21.360000 128.135000 23.160000 129.385000 ;
        RECT 21.360000 119.995000 23.160000 121.245000 ;
        RECT 10.560000 152.555000 12.360000 153.805000 ;
        RECT 10.560000 144.415000 12.360000 145.665000 ;
        RECT 7.360000 144.415000 9.360000 145.665000 ;
        RECT 7.360000 152.555000 9.360000 153.805000 ;
        RECT 32.160000 152.555000 33.960000 153.805000 ;
        RECT 32.160000 144.415000 33.960000 145.665000 ;
        RECT 21.360000 152.555000 23.160000 153.805000 ;
        RECT 21.360000 144.415000 23.160000 145.665000 ;
        RECT 75.360000 136.275000 77.160000 137.525000 ;
        RECT 64.560000 136.275000 66.360000 137.525000 ;
        RECT 53.760000 136.275000 55.560000 137.525000 ;
        RECT 42.960000 136.275000 44.760000 137.525000 ;
        RECT 42.960000 119.995000 44.760000 121.245000 ;
        RECT 42.960000 128.135000 44.760000 129.385000 ;
        RECT 53.760000 119.995000 55.560000 121.245000 ;
        RECT 53.760000 128.135000 55.560000 129.385000 ;
        RECT 64.560000 119.995000 66.360000 121.245000 ;
        RECT 64.560000 128.135000 66.360000 129.385000 ;
        RECT 75.360000 119.995000 77.160000 121.245000 ;
        RECT 75.360000 128.135000 77.160000 129.385000 ;
        RECT 42.960000 144.415000 44.760000 145.665000 ;
        RECT 42.960000 152.555000 44.760000 153.805000 ;
        RECT 53.760000 144.415000 55.560000 145.665000 ;
        RECT 53.760000 152.555000 55.560000 153.805000 ;
        RECT 64.560000 144.415000 66.360000 145.665000 ;
        RECT 64.560000 152.555000 66.360000 153.805000 ;
        RECT 75.360000 144.415000 77.160000 145.665000 ;
        RECT 75.360000 152.555000 77.160000 153.805000 ;
        RECT 96.960000 95.575000 98.760000 96.825000 ;
        RECT 96.960000 87.435000 98.760000 88.685000 ;
        RECT 96.960000 79.295000 98.760000 80.545000 ;
        RECT 86.160000 79.295000 87.960000 80.545000 ;
        RECT 86.160000 87.435000 87.960000 88.685000 ;
        RECT 86.160000 95.575000 87.960000 96.825000 ;
        RECT 107.760000 95.575000 109.560000 96.825000 ;
        RECT 107.760000 87.435000 109.560000 88.685000 ;
        RECT 107.760000 79.295000 109.560000 80.545000 ;
        RECT 96.960000 111.855000 98.760000 113.105000 ;
        RECT 96.960000 103.715000 98.760000 104.965000 ;
        RECT 86.160000 103.715000 87.960000 104.965000 ;
        RECT 86.160000 111.855000 87.960000 113.105000 ;
        RECT 107.760000 103.715000 109.560000 104.965000 ;
        RECT 107.760000 111.855000 109.560000 113.105000 ;
        RECT 118.560000 87.435000 120.360000 88.685000 ;
        RECT 129.360000 87.435000 131.160000 88.685000 ;
        RECT 129.360000 79.295000 131.160000 80.545000 ;
        RECT 118.560000 79.295000 120.360000 80.545000 ;
        RECT 129.360000 95.575000 131.160000 96.825000 ;
        RECT 118.560000 95.575000 120.360000 96.825000 ;
        RECT 140.160000 79.295000 141.960000 80.545000 ;
        RECT 140.160000 87.435000 141.960000 88.685000 ;
        RECT 140.160000 95.575000 141.960000 96.825000 ;
        RECT 150.960000 79.295000 152.760000 80.545000 ;
        RECT 150.960000 87.435000 152.760000 88.685000 ;
        RECT 150.960000 95.575000 152.760000 96.825000 ;
        RECT 118.560000 103.715000 120.360000 104.965000 ;
        RECT 118.560000 111.855000 120.360000 113.105000 ;
        RECT 129.360000 103.715000 131.160000 104.965000 ;
        RECT 129.360000 111.855000 131.160000 113.105000 ;
        RECT 140.160000 103.715000 141.960000 104.965000 ;
        RECT 140.160000 111.855000 141.960000 113.105000 ;
        RECT 150.960000 103.715000 152.760000 104.965000 ;
        RECT 150.960000 111.855000 152.760000 113.105000 ;
        RECT 107.760000 136.275000 109.560000 137.525000 ;
        RECT 96.960000 136.275000 98.760000 137.525000 ;
        RECT 86.160000 136.275000 87.960000 137.525000 ;
        RECT 96.960000 128.135000 98.760000 129.385000 ;
        RECT 96.960000 119.995000 98.760000 121.245000 ;
        RECT 86.160000 119.995000 87.960000 121.245000 ;
        RECT 86.160000 128.135000 87.960000 129.385000 ;
        RECT 107.760000 119.995000 109.560000 121.245000 ;
        RECT 107.760000 128.135000 109.560000 129.385000 ;
        RECT 96.960000 152.555000 98.760000 153.805000 ;
        RECT 96.960000 144.415000 98.760000 145.665000 ;
        RECT 86.160000 144.415000 87.960000 145.665000 ;
        RECT 86.160000 152.555000 87.960000 153.805000 ;
        RECT 107.760000 144.415000 109.560000 145.665000 ;
        RECT 107.760000 152.555000 109.560000 153.805000 ;
        RECT 150.960000 136.275000 152.760000 137.525000 ;
        RECT 140.160000 136.275000 141.960000 137.525000 ;
        RECT 129.360000 136.275000 131.160000 137.525000 ;
        RECT 118.560000 136.275000 120.360000 137.525000 ;
        RECT 118.560000 119.995000 120.360000 121.245000 ;
        RECT 118.560000 128.135000 120.360000 129.385000 ;
        RECT 129.360000 119.995000 131.160000 121.245000 ;
        RECT 129.360000 128.135000 131.160000 129.385000 ;
        RECT 140.160000 119.995000 141.960000 121.245000 ;
        RECT 140.160000 128.135000 141.960000 129.385000 ;
        RECT 150.960000 119.995000 152.760000 121.245000 ;
        RECT 150.960000 128.135000 152.760000 129.385000 ;
        RECT 118.560000 144.415000 120.360000 145.665000 ;
        RECT 118.560000 152.555000 120.360000 153.805000 ;
        RECT 129.360000 144.415000 131.160000 145.665000 ;
        RECT 129.360000 152.555000 131.160000 153.805000 ;
        RECT 140.160000 144.415000 141.960000 145.665000 ;
        RECT 140.160000 152.555000 141.960000 153.805000 ;
        RECT 150.960000 144.415000 152.760000 145.665000 ;
        RECT 150.960000 152.555000 152.760000 153.805000 ;
        RECT 226.560000 38.595000 228.360000 39.845000 ;
        RECT 215.760000 38.595000 217.560000 39.845000 ;
        RECT 204.960000 38.595000 206.760000 39.845000 ;
        RECT 194.160000 38.595000 195.960000 39.845000 ;
        RECT 183.360000 38.595000 185.160000 39.845000 ;
        RECT 172.560000 38.595000 174.360000 39.845000 ;
        RECT 161.760000 38.595000 163.560000 39.845000 ;
        RECT 194.160000 30.455000 195.960000 31.705000 ;
        RECT 194.160000 22.315000 195.960000 23.565000 ;
        RECT 194.160000 14.175000 195.960000 15.425000 ;
        RECT 183.360000 14.175000 185.160000 15.425000 ;
        RECT 172.560000 14.175000 174.360000 15.425000 ;
        RECT 161.760000 14.175000 163.560000 15.425000 ;
        RECT 183.360000 30.455000 185.160000 31.705000 ;
        RECT 183.360000 22.315000 185.160000 23.565000 ;
        RECT 172.560000 30.455000 174.360000 31.705000 ;
        RECT 172.560000 22.315000 174.360000 23.565000 ;
        RECT 161.760000 30.455000 163.560000 31.705000 ;
        RECT 161.760000 22.315000 163.560000 23.565000 ;
        RECT 215.760000 14.175000 217.560000 15.425000 ;
        RECT 204.960000 14.175000 206.760000 15.425000 ;
        RECT 226.560000 14.175000 228.360000 15.425000 ;
        RECT 204.960000 30.455000 206.760000 31.705000 ;
        RECT 204.960000 22.315000 206.760000 23.565000 ;
        RECT 215.760000 22.315000 217.560000 23.565000 ;
        RECT 215.760000 30.455000 217.560000 31.705000 ;
        RECT 226.560000 22.315000 228.360000 23.565000 ;
        RECT 226.560000 30.455000 228.360000 31.705000 ;
        RECT 194.160000 71.155000 195.960000 72.405000 ;
        RECT 194.160000 63.015000 195.960000 64.265000 ;
        RECT 194.160000 54.875000 195.960000 56.125000 ;
        RECT 194.160000 46.735000 195.960000 47.985000 ;
        RECT 183.360000 46.735000 185.160000 47.985000 ;
        RECT 172.560000 54.875000 174.360000 56.125000 ;
        RECT 172.560000 46.735000 174.360000 47.985000 ;
        RECT 161.760000 54.875000 163.560000 56.125000 ;
        RECT 161.760000 46.735000 163.560000 47.985000 ;
        RECT 183.360000 54.875000 185.160000 56.125000 ;
        RECT 172.560000 71.155000 174.360000 72.405000 ;
        RECT 172.560000 63.015000 174.360000 64.265000 ;
        RECT 161.760000 71.155000 163.560000 72.405000 ;
        RECT 161.760000 63.015000 163.560000 64.265000 ;
        RECT 183.360000 63.015000 185.160000 64.265000 ;
        RECT 183.360000 71.155000 185.160000 72.405000 ;
        RECT 204.960000 46.735000 206.760000 47.985000 ;
        RECT 204.960000 54.875000 206.760000 56.125000 ;
        RECT 215.760000 46.735000 217.560000 47.985000 ;
        RECT 215.760000 54.875000 217.560000 56.125000 ;
        RECT 226.560000 46.735000 228.360000 47.985000 ;
        RECT 226.560000 54.875000 228.360000 56.125000 ;
        RECT 204.960000 71.155000 206.760000 72.405000 ;
        RECT 204.960000 63.015000 206.760000 64.265000 ;
        RECT 226.560000 71.155000 228.360000 72.405000 ;
        RECT 226.560000 63.015000 228.360000 64.265000 ;
        RECT 215.760000 71.155000 217.560000 72.405000 ;
        RECT 215.760000 63.015000 217.560000 64.265000 ;
        RECT 291.360000 38.595000 293.160000 39.845000 ;
        RECT 280.560000 38.595000 282.360000 39.845000 ;
        RECT 269.760000 38.595000 271.560000 39.845000 ;
        RECT 258.960000 38.595000 260.760000 39.845000 ;
        RECT 248.160000 38.595000 249.960000 39.845000 ;
        RECT 237.360000 38.595000 239.160000 39.845000 ;
        RECT 301.680000 38.595000 303.680000 39.845000 ;
        RECT 237.360000 14.175000 239.160000 15.425000 ;
        RECT 248.160000 14.175000 249.960000 15.425000 ;
        RECT 258.960000 14.175000 260.760000 15.425000 ;
        RECT 269.760000 14.175000 271.560000 15.425000 ;
        RECT 237.360000 22.315000 239.160000 23.565000 ;
        RECT 237.360000 30.455000 239.160000 31.705000 ;
        RECT 248.160000 22.315000 249.960000 23.565000 ;
        RECT 248.160000 30.455000 249.960000 31.705000 ;
        RECT 258.960000 22.315000 260.760000 23.565000 ;
        RECT 258.960000 30.455000 260.760000 31.705000 ;
        RECT 269.760000 22.315000 271.560000 23.565000 ;
        RECT 269.760000 30.455000 271.560000 31.705000 ;
        RECT 291.360000 14.175000 293.160000 15.425000 ;
        RECT 301.680000 14.175000 303.680000 15.425000 ;
        RECT 280.560000 14.175000 282.360000 15.425000 ;
        RECT 291.360000 30.455000 293.160000 31.705000 ;
        RECT 291.360000 22.315000 293.160000 23.565000 ;
        RECT 280.560000 30.455000 282.360000 31.705000 ;
        RECT 280.560000 22.315000 282.360000 23.565000 ;
        RECT 301.680000 30.455000 303.680000 31.705000 ;
        RECT 301.680000 22.315000 303.680000 23.565000 ;
        RECT 237.360000 46.735000 239.160000 47.985000 ;
        RECT 237.360000 54.875000 239.160000 56.125000 ;
        RECT 248.160000 46.735000 249.960000 47.985000 ;
        RECT 248.160000 54.875000 249.960000 56.125000 ;
        RECT 258.960000 46.735000 260.760000 47.985000 ;
        RECT 258.960000 54.875000 260.760000 56.125000 ;
        RECT 269.760000 46.735000 271.560000 47.985000 ;
        RECT 269.760000 54.875000 271.560000 56.125000 ;
        RECT 248.160000 71.155000 249.960000 72.405000 ;
        RECT 248.160000 63.015000 249.960000 64.265000 ;
        RECT 237.360000 71.155000 239.160000 72.405000 ;
        RECT 237.360000 63.015000 239.160000 64.265000 ;
        RECT 269.760000 71.155000 271.560000 72.405000 ;
        RECT 269.760000 63.015000 271.560000 64.265000 ;
        RECT 258.960000 71.155000 260.760000 72.405000 ;
        RECT 258.960000 63.015000 260.760000 64.265000 ;
        RECT 291.360000 54.875000 293.160000 56.125000 ;
        RECT 291.360000 46.735000 293.160000 47.985000 ;
        RECT 280.560000 54.875000 282.360000 56.125000 ;
        RECT 280.560000 46.735000 282.360000 47.985000 ;
        RECT 301.680000 54.875000 303.680000 56.125000 ;
        RECT 301.680000 46.735000 303.680000 47.985000 ;
        RECT 291.360000 71.155000 293.160000 72.405000 ;
        RECT 291.360000 63.015000 293.160000 64.265000 ;
        RECT 280.560000 63.015000 282.360000 64.265000 ;
        RECT 280.560000 71.155000 282.360000 72.405000 ;
        RECT 301.680000 63.015000 303.680000 64.265000 ;
        RECT 301.680000 71.155000 303.680000 72.405000 ;
        RECT 194.160000 111.855000 195.960000 113.105000 ;
        RECT 194.160000 103.715000 195.960000 104.965000 ;
        RECT 194.160000 95.575000 195.960000 96.825000 ;
        RECT 194.160000 87.435000 195.960000 88.685000 ;
        RECT 194.160000 79.295000 195.960000 80.545000 ;
        RECT 161.760000 79.295000 163.560000 80.545000 ;
        RECT 161.760000 87.435000 163.560000 88.685000 ;
        RECT 161.760000 95.575000 163.560000 96.825000 ;
        RECT 172.560000 79.295000 174.360000 80.545000 ;
        RECT 172.560000 87.435000 174.360000 88.685000 ;
        RECT 172.560000 95.575000 174.360000 96.825000 ;
        RECT 183.360000 79.295000 185.160000 80.545000 ;
        RECT 183.360000 87.435000 185.160000 88.685000 ;
        RECT 183.360000 95.575000 185.160000 96.825000 ;
        RECT 161.760000 103.715000 163.560000 104.965000 ;
        RECT 161.760000 111.855000 163.560000 113.105000 ;
        RECT 172.560000 103.715000 174.360000 104.965000 ;
        RECT 172.560000 111.855000 174.360000 113.105000 ;
        RECT 183.360000 103.715000 185.160000 104.965000 ;
        RECT 183.360000 111.855000 185.160000 113.105000 ;
        RECT 204.960000 79.295000 206.760000 80.545000 ;
        RECT 204.960000 87.435000 206.760000 88.685000 ;
        RECT 204.960000 95.575000 206.760000 96.825000 ;
        RECT 226.560000 87.435000 228.360000 88.685000 ;
        RECT 215.760000 87.435000 217.560000 88.685000 ;
        RECT 215.760000 79.295000 217.560000 80.545000 ;
        RECT 226.560000 79.295000 228.360000 80.545000 ;
        RECT 215.760000 95.575000 217.560000 96.825000 ;
        RECT 226.560000 95.575000 228.360000 96.825000 ;
        RECT 204.960000 103.715000 206.760000 104.965000 ;
        RECT 204.960000 111.855000 206.760000 113.105000 ;
        RECT 215.760000 103.715000 217.560000 104.965000 ;
        RECT 215.760000 111.855000 217.560000 113.105000 ;
        RECT 226.560000 103.715000 228.360000 104.965000 ;
        RECT 226.560000 111.855000 228.360000 113.105000 ;
        RECT 194.160000 152.555000 195.960000 153.805000 ;
        RECT 194.160000 144.415000 195.960000 145.665000 ;
        RECT 194.160000 136.275000 195.960000 137.525000 ;
        RECT 194.160000 128.135000 195.960000 129.385000 ;
        RECT 194.160000 119.995000 195.960000 121.245000 ;
        RECT 183.360000 136.275000 185.160000 137.525000 ;
        RECT 172.560000 136.275000 174.360000 137.525000 ;
        RECT 161.760000 136.275000 163.560000 137.525000 ;
        RECT 161.760000 119.995000 163.560000 121.245000 ;
        RECT 161.760000 128.135000 163.560000 129.385000 ;
        RECT 172.560000 119.995000 174.360000 121.245000 ;
        RECT 172.560000 128.135000 174.360000 129.385000 ;
        RECT 183.360000 119.995000 185.160000 121.245000 ;
        RECT 183.360000 128.135000 185.160000 129.385000 ;
        RECT 161.760000 144.415000 163.560000 145.665000 ;
        RECT 161.760000 152.555000 163.560000 153.805000 ;
        RECT 172.560000 144.415000 174.360000 145.665000 ;
        RECT 172.560000 152.555000 174.360000 153.805000 ;
        RECT 183.360000 144.415000 185.160000 145.665000 ;
        RECT 183.360000 152.555000 185.160000 153.805000 ;
        RECT 226.560000 136.275000 228.360000 137.525000 ;
        RECT 215.760000 136.275000 217.560000 137.525000 ;
        RECT 204.960000 136.275000 206.760000 137.525000 ;
        RECT 204.960000 119.995000 206.760000 121.245000 ;
        RECT 204.960000 128.135000 206.760000 129.385000 ;
        RECT 215.760000 119.995000 217.560000 121.245000 ;
        RECT 215.760000 128.135000 217.560000 129.385000 ;
        RECT 226.560000 119.995000 228.360000 121.245000 ;
        RECT 226.560000 128.135000 228.360000 129.385000 ;
        RECT 204.960000 144.415000 206.760000 145.665000 ;
        RECT 204.960000 152.555000 206.760000 153.805000 ;
        RECT 215.760000 144.415000 217.560000 145.665000 ;
        RECT 215.760000 152.555000 217.560000 153.805000 ;
        RECT 226.560000 144.415000 228.360000 145.665000 ;
        RECT 226.560000 152.555000 228.360000 153.805000 ;
        RECT 237.360000 79.295000 239.160000 80.545000 ;
        RECT 237.360000 87.435000 239.160000 88.685000 ;
        RECT 237.360000 95.575000 239.160000 96.825000 ;
        RECT 248.160000 79.295000 249.960000 80.545000 ;
        RECT 248.160000 87.435000 249.960000 88.685000 ;
        RECT 248.160000 95.575000 249.960000 96.825000 ;
        RECT 258.960000 79.295000 260.760000 80.545000 ;
        RECT 258.960000 87.435000 260.760000 88.685000 ;
        RECT 258.960000 95.575000 260.760000 96.825000 ;
        RECT 269.760000 79.295000 271.560000 80.545000 ;
        RECT 269.760000 87.435000 271.560000 88.685000 ;
        RECT 269.760000 95.575000 271.560000 96.825000 ;
        RECT 237.360000 103.715000 239.160000 104.965000 ;
        RECT 237.360000 111.855000 239.160000 113.105000 ;
        RECT 248.160000 103.715000 249.960000 104.965000 ;
        RECT 248.160000 111.855000 249.960000 113.105000 ;
        RECT 258.960000 103.715000 260.760000 104.965000 ;
        RECT 258.960000 111.855000 260.760000 113.105000 ;
        RECT 269.760000 103.715000 271.560000 104.965000 ;
        RECT 269.760000 111.855000 271.560000 113.105000 ;
        RECT 291.360000 95.575000 293.160000 96.825000 ;
        RECT 291.360000 87.435000 293.160000 88.685000 ;
        RECT 291.360000 79.295000 293.160000 80.545000 ;
        RECT 280.560000 95.575000 282.360000 96.825000 ;
        RECT 280.560000 87.435000 282.360000 88.685000 ;
        RECT 280.560000 79.295000 282.360000 80.545000 ;
        RECT 301.680000 95.575000 303.680000 96.825000 ;
        RECT 301.680000 87.435000 303.680000 88.685000 ;
        RECT 301.680000 79.295000 303.680000 80.545000 ;
        RECT 291.360000 111.855000 293.160000 113.105000 ;
        RECT 291.360000 103.715000 293.160000 104.965000 ;
        RECT 280.560000 111.855000 282.360000 113.105000 ;
        RECT 280.560000 103.715000 282.360000 104.965000 ;
        RECT 301.680000 103.715000 303.680000 104.965000 ;
        RECT 301.680000 111.855000 303.680000 113.105000 ;
        RECT 269.760000 136.275000 271.560000 137.525000 ;
        RECT 258.960000 136.275000 260.760000 137.525000 ;
        RECT 248.160000 136.275000 249.960000 137.525000 ;
        RECT 237.360000 136.275000 239.160000 137.525000 ;
        RECT 237.360000 119.995000 239.160000 121.245000 ;
        RECT 237.360000 128.135000 239.160000 129.385000 ;
        RECT 248.160000 119.995000 249.960000 121.245000 ;
        RECT 248.160000 128.135000 249.960000 129.385000 ;
        RECT 258.960000 119.995000 260.760000 121.245000 ;
        RECT 258.960000 128.135000 260.760000 129.385000 ;
        RECT 269.760000 119.995000 271.560000 121.245000 ;
        RECT 269.760000 128.135000 271.560000 129.385000 ;
        RECT 237.360000 144.415000 239.160000 145.665000 ;
        RECT 237.360000 152.555000 239.160000 153.805000 ;
        RECT 248.160000 144.415000 249.960000 145.665000 ;
        RECT 248.160000 152.555000 249.960000 153.805000 ;
        RECT 258.960000 144.415000 260.760000 145.665000 ;
        RECT 258.960000 152.555000 260.760000 153.805000 ;
        RECT 269.760000 144.415000 271.560000 145.665000 ;
        RECT 269.760000 152.555000 271.560000 153.805000 ;
        RECT 291.360000 136.275000 293.160000 137.525000 ;
        RECT 280.560000 136.275000 282.360000 137.525000 ;
        RECT 301.680000 136.275000 303.680000 137.525000 ;
        RECT 291.360000 128.135000 293.160000 129.385000 ;
        RECT 291.360000 119.995000 293.160000 121.245000 ;
        RECT 280.560000 128.135000 282.360000 129.385000 ;
        RECT 280.560000 119.995000 282.360000 121.245000 ;
        RECT 301.680000 119.995000 303.680000 121.245000 ;
        RECT 301.680000 128.135000 303.680000 129.385000 ;
        RECT 291.360000 152.555000 293.160000 153.805000 ;
        RECT 291.360000 144.415000 293.160000 145.665000 ;
        RECT 280.560000 152.555000 282.360000 153.805000 ;
        RECT 280.560000 144.415000 282.360000 145.665000 ;
        RECT 301.680000 144.415000 303.680000 145.665000 ;
        RECT 301.680000 152.555000 303.680000 153.805000 ;
        RECT 7.360000 160.695000 9.360000 161.945000 ;
        RECT 10.560000 160.695000 12.360000 161.945000 ;
        RECT 7.360000 168.835000 9.360000 170.085000 ;
        RECT 10.560000 168.835000 12.360000 170.085000 ;
        RECT 21.360000 160.695000 23.160000 161.945000 ;
        RECT 32.160000 160.695000 33.960000 161.945000 ;
        RECT 21.360000 168.835000 23.160000 170.085000 ;
        RECT 32.160000 168.835000 33.960000 170.085000 ;
        RECT 7.360000 176.975000 9.360000 178.225000 ;
        RECT 10.560000 176.975000 12.360000 178.225000 ;
        RECT 7.360000 185.115000 9.360000 186.365000 ;
        RECT 7.360000 193.255000 9.360000 194.505000 ;
        RECT 10.560000 185.115000 12.360000 186.365000 ;
        RECT 10.560000 193.255000 12.360000 194.505000 ;
        RECT 21.360000 176.975000 23.160000 178.225000 ;
        RECT 32.160000 176.975000 33.960000 178.225000 ;
        RECT 21.360000 185.115000 23.160000 186.365000 ;
        RECT 21.360000 193.255000 23.160000 194.505000 ;
        RECT 32.160000 185.115000 33.960000 186.365000 ;
        RECT 32.160000 193.255000 33.960000 194.505000 ;
        RECT 53.760000 168.835000 55.560000 170.085000 ;
        RECT 42.960000 160.695000 44.760000 161.945000 ;
        RECT 42.960000 168.835000 44.760000 170.085000 ;
        RECT 53.760000 160.695000 55.560000 161.945000 ;
        RECT 75.360000 168.835000 77.160000 170.085000 ;
        RECT 75.360000 160.695000 77.160000 161.945000 ;
        RECT 64.560000 168.835000 66.360000 170.085000 ;
        RECT 64.560000 160.695000 66.360000 161.945000 ;
        RECT 42.960000 176.975000 44.760000 178.225000 ;
        RECT 42.960000 185.115000 44.760000 186.365000 ;
        RECT 42.960000 193.255000 44.760000 194.505000 ;
        RECT 53.760000 176.975000 55.560000 178.225000 ;
        RECT 53.760000 185.115000 55.560000 186.365000 ;
        RECT 53.760000 193.255000 55.560000 194.505000 ;
        RECT 64.560000 176.975000 66.360000 178.225000 ;
        RECT 64.560000 185.115000 66.360000 186.365000 ;
        RECT 64.560000 193.255000 66.360000 194.505000 ;
        RECT 75.360000 176.975000 77.160000 178.225000 ;
        RECT 75.360000 185.115000 77.160000 186.365000 ;
        RECT 75.360000 193.255000 77.160000 194.505000 ;
        RECT 10.560000 209.535000 12.360000 210.785000 ;
        RECT 10.560000 201.395000 12.360000 202.645000 ;
        RECT 7.360000 201.395000 9.360000 202.645000 ;
        RECT 7.360000 209.535000 9.360000 210.785000 ;
        RECT 32.160000 209.535000 33.960000 210.785000 ;
        RECT 32.160000 201.395000 33.960000 202.645000 ;
        RECT 21.360000 209.535000 23.160000 210.785000 ;
        RECT 21.360000 201.395000 23.160000 202.645000 ;
        RECT 10.560000 225.815000 12.360000 227.065000 ;
        RECT 10.560000 217.675000 12.360000 218.925000 ;
        RECT 7.360000 217.675000 9.360000 218.925000 ;
        RECT 7.360000 225.815000 9.360000 227.065000 ;
        RECT 32.160000 225.815000 33.960000 227.065000 ;
        RECT 32.160000 217.675000 33.960000 218.925000 ;
        RECT 21.360000 225.815000 23.160000 227.065000 ;
        RECT 21.360000 217.675000 23.160000 218.925000 ;
        RECT 42.960000 201.395000 44.760000 202.645000 ;
        RECT 42.960000 209.535000 44.760000 210.785000 ;
        RECT 53.760000 201.395000 55.560000 202.645000 ;
        RECT 53.760000 209.535000 55.560000 210.785000 ;
        RECT 64.560000 201.395000 66.360000 202.645000 ;
        RECT 64.560000 209.535000 66.360000 210.785000 ;
        RECT 75.360000 201.395000 77.160000 202.645000 ;
        RECT 75.360000 209.535000 77.160000 210.785000 ;
        RECT 42.960000 217.675000 44.760000 218.925000 ;
        RECT 42.960000 225.815000 44.760000 227.065000 ;
        RECT 53.760000 217.675000 55.560000 218.925000 ;
        RECT 53.760000 225.815000 55.560000 227.065000 ;
        RECT 64.560000 217.675000 66.360000 218.925000 ;
        RECT 64.560000 225.815000 66.360000 227.065000 ;
        RECT 75.360000 217.675000 77.160000 218.925000 ;
        RECT 75.360000 225.815000 77.160000 227.065000 ;
        RECT 96.960000 168.835000 98.760000 170.085000 ;
        RECT 96.960000 160.695000 98.760000 161.945000 ;
        RECT 86.160000 168.835000 87.960000 170.085000 ;
        RECT 86.160000 160.695000 87.960000 161.945000 ;
        RECT 107.760000 168.835000 109.560000 170.085000 ;
        RECT 107.760000 160.695000 109.560000 161.945000 ;
        RECT 96.960000 193.255000 98.760000 194.505000 ;
        RECT 96.960000 185.115000 98.760000 186.365000 ;
        RECT 96.960000 176.975000 98.760000 178.225000 ;
        RECT 86.160000 176.975000 87.960000 178.225000 ;
        RECT 86.160000 185.115000 87.960000 186.365000 ;
        RECT 86.160000 193.255000 87.960000 194.505000 ;
        RECT 107.760000 193.255000 109.560000 194.505000 ;
        RECT 107.760000 185.115000 109.560000 186.365000 ;
        RECT 107.760000 176.975000 109.560000 178.225000 ;
        RECT 129.360000 160.695000 131.160000 161.945000 ;
        RECT 118.560000 160.695000 120.360000 161.945000 ;
        RECT 118.560000 168.835000 120.360000 170.085000 ;
        RECT 129.360000 168.835000 131.160000 170.085000 ;
        RECT 150.960000 168.835000 152.760000 170.085000 ;
        RECT 150.960000 160.695000 152.760000 161.945000 ;
        RECT 140.160000 168.835000 141.960000 170.085000 ;
        RECT 140.160000 160.695000 141.960000 161.945000 ;
        RECT 129.360000 176.975000 131.160000 178.225000 ;
        RECT 118.560000 176.975000 120.360000 178.225000 ;
        RECT 129.360000 193.255000 131.160000 194.505000 ;
        RECT 129.360000 185.115000 131.160000 186.365000 ;
        RECT 118.560000 193.255000 120.360000 194.505000 ;
        RECT 118.560000 185.115000 120.360000 186.365000 ;
        RECT 140.160000 176.975000 141.960000 178.225000 ;
        RECT 140.160000 185.115000 141.960000 186.365000 ;
        RECT 140.160000 193.255000 141.960000 194.505000 ;
        RECT 150.960000 176.975000 152.760000 178.225000 ;
        RECT 150.960000 185.115000 152.760000 186.365000 ;
        RECT 150.960000 193.255000 152.760000 194.505000 ;
        RECT 96.960000 209.535000 98.760000 210.785000 ;
        RECT 96.960000 201.395000 98.760000 202.645000 ;
        RECT 86.160000 201.395000 87.960000 202.645000 ;
        RECT 86.160000 209.535000 87.960000 210.785000 ;
        RECT 107.760000 201.395000 109.560000 202.645000 ;
        RECT 107.760000 209.535000 109.560000 210.785000 ;
        RECT 96.960000 225.815000 98.760000 227.065000 ;
        RECT 96.960000 217.675000 98.760000 218.925000 ;
        RECT 86.160000 217.675000 87.960000 218.925000 ;
        RECT 86.160000 225.815000 87.960000 227.065000 ;
        RECT 107.760000 217.675000 109.560000 218.925000 ;
        RECT 107.760000 225.815000 109.560000 227.065000 ;
        RECT 118.560000 201.395000 120.360000 202.645000 ;
        RECT 118.560000 209.535000 120.360000 210.785000 ;
        RECT 129.360000 201.395000 131.160000 202.645000 ;
        RECT 129.360000 209.535000 131.160000 210.785000 ;
        RECT 140.160000 201.395000 141.960000 202.645000 ;
        RECT 140.160000 209.535000 141.960000 210.785000 ;
        RECT 150.960000 201.395000 152.760000 202.645000 ;
        RECT 150.960000 209.535000 152.760000 210.785000 ;
        RECT 118.560000 217.675000 120.360000 218.925000 ;
        RECT 118.560000 225.815000 120.360000 227.065000 ;
        RECT 129.360000 217.675000 131.160000 218.925000 ;
        RECT 129.360000 225.815000 131.160000 227.065000 ;
        RECT 140.160000 217.675000 141.960000 218.925000 ;
        RECT 140.160000 225.815000 141.960000 227.065000 ;
        RECT 150.960000 217.675000 152.760000 218.925000 ;
        RECT 150.960000 225.815000 152.760000 227.065000 ;
        RECT 7.360000 233.955000 9.360000 235.205000 ;
        RECT 7.360000 242.095000 9.360000 243.345000 ;
        RECT 10.560000 233.955000 12.360000 235.205000 ;
        RECT 10.560000 242.095000 12.360000 243.345000 ;
        RECT 7.360000 250.235000 9.360000 251.485000 ;
        RECT 10.560000 250.235000 12.360000 251.485000 ;
        RECT 21.360000 233.955000 23.160000 235.205000 ;
        RECT 21.360000 242.095000 23.160000 243.345000 ;
        RECT 32.160000 233.955000 33.960000 235.205000 ;
        RECT 32.160000 242.095000 33.960000 243.345000 ;
        RECT 21.360000 250.235000 23.160000 251.485000 ;
        RECT 32.160000 250.235000 33.960000 251.485000 ;
        RECT 7.360000 258.375000 9.360000 259.625000 ;
        RECT 10.560000 258.375000 12.360000 259.625000 ;
        RECT 7.360000 266.515000 9.360000 267.765000 ;
        RECT 10.560000 266.515000 12.360000 267.765000 ;
        RECT 21.360000 258.375000 23.160000 259.625000 ;
        RECT 32.160000 258.375000 33.960000 259.625000 ;
        RECT 21.360000 266.515000 23.160000 267.765000 ;
        RECT 32.160000 266.515000 33.960000 267.765000 ;
        RECT 42.960000 233.955000 44.760000 235.205000 ;
        RECT 42.960000 242.095000 44.760000 243.345000 ;
        RECT 42.960000 250.235000 44.760000 251.485000 ;
        RECT 53.760000 233.955000 55.560000 235.205000 ;
        RECT 53.760000 242.095000 55.560000 243.345000 ;
        RECT 53.760000 250.235000 55.560000 251.485000 ;
        RECT 64.560000 233.955000 66.360000 235.205000 ;
        RECT 64.560000 242.095000 66.360000 243.345000 ;
        RECT 64.560000 250.235000 66.360000 251.485000 ;
        RECT 75.360000 233.955000 77.160000 235.205000 ;
        RECT 75.360000 242.095000 77.160000 243.345000 ;
        RECT 75.360000 250.235000 77.160000 251.485000 ;
        RECT 53.760000 266.515000 55.560000 267.765000 ;
        RECT 42.960000 258.375000 44.760000 259.625000 ;
        RECT 42.960000 266.515000 44.760000 267.765000 ;
        RECT 53.760000 258.375000 55.560000 259.625000 ;
        RECT 75.360000 266.515000 77.160000 267.765000 ;
        RECT 75.360000 258.375000 77.160000 259.625000 ;
        RECT 64.560000 266.515000 66.360000 267.765000 ;
        RECT 64.560000 258.375000 66.360000 259.625000 ;
        RECT 32.160000 290.935000 33.960000 292.185000 ;
        RECT 21.360000 290.935000 23.160000 292.185000 ;
        RECT 10.560000 290.935000 12.360000 292.185000 ;
        RECT 7.360000 290.935000 9.360000 292.185000 ;
        RECT 10.560000 282.795000 12.360000 284.045000 ;
        RECT 10.560000 274.655000 12.360000 275.905000 ;
        RECT 7.360000 274.655000 9.360000 275.905000 ;
        RECT 7.360000 282.795000 9.360000 284.045000 ;
        RECT 32.160000 282.795000 33.960000 284.045000 ;
        RECT 32.160000 274.655000 33.960000 275.905000 ;
        RECT 21.360000 282.795000 23.160000 284.045000 ;
        RECT 21.360000 274.655000 23.160000 275.905000 ;
        RECT 9.785000 298.940000 10.165000 299.580000 ;
        RECT 7.360000 299.535000 9.360000 299.865000 ;
        RECT 10.560000 299.075000 12.360000 299.865000 ;
        RECT 32.160000 299.075000 33.960000 299.865000 ;
        RECT 21.360000 299.075000 23.160000 299.865000 ;
        RECT 75.360000 290.935000 77.160000 292.185000 ;
        RECT 64.560000 290.935000 66.360000 292.185000 ;
        RECT 53.760000 290.935000 55.560000 292.185000 ;
        RECT 42.960000 290.935000 44.760000 292.185000 ;
        RECT 42.960000 274.655000 44.760000 275.905000 ;
        RECT 42.960000 282.795000 44.760000 284.045000 ;
        RECT 53.760000 274.655000 55.560000 275.905000 ;
        RECT 53.760000 282.795000 55.560000 284.045000 ;
        RECT 64.560000 274.655000 66.360000 275.905000 ;
        RECT 64.560000 282.795000 66.360000 284.045000 ;
        RECT 75.360000 274.655000 77.160000 275.905000 ;
        RECT 75.360000 282.795000 77.160000 284.045000 ;
        RECT 42.960000 299.075000 44.760000 299.865000 ;
        RECT 53.760000 299.075000 55.560000 299.865000 ;
        RECT 64.560000 299.075000 66.360000 299.865000 ;
        RECT 75.360000 299.075000 77.160000 299.865000 ;
        RECT 96.960000 250.235000 98.760000 251.485000 ;
        RECT 96.960000 242.095000 98.760000 243.345000 ;
        RECT 96.960000 233.955000 98.760000 235.205000 ;
        RECT 86.160000 233.955000 87.960000 235.205000 ;
        RECT 86.160000 242.095000 87.960000 243.345000 ;
        RECT 86.160000 250.235000 87.960000 251.485000 ;
        RECT 107.760000 250.235000 109.560000 251.485000 ;
        RECT 107.760000 242.095000 109.560000 243.345000 ;
        RECT 107.760000 233.955000 109.560000 235.205000 ;
        RECT 96.960000 266.515000 98.760000 267.765000 ;
        RECT 96.960000 258.375000 98.760000 259.625000 ;
        RECT 86.160000 266.515000 87.960000 267.765000 ;
        RECT 86.160000 258.375000 87.960000 259.625000 ;
        RECT 107.760000 266.515000 109.560000 267.765000 ;
        RECT 107.760000 258.375000 109.560000 259.625000 ;
        RECT 129.360000 242.095000 131.160000 243.345000 ;
        RECT 129.360000 233.955000 131.160000 235.205000 ;
        RECT 118.560000 242.095000 120.360000 243.345000 ;
        RECT 118.560000 233.955000 120.360000 235.205000 ;
        RECT 129.360000 250.235000 131.160000 251.485000 ;
        RECT 118.560000 250.235000 120.360000 251.485000 ;
        RECT 140.160000 233.955000 141.960000 235.205000 ;
        RECT 140.160000 242.095000 141.960000 243.345000 ;
        RECT 140.160000 250.235000 141.960000 251.485000 ;
        RECT 150.960000 233.955000 152.760000 235.205000 ;
        RECT 150.960000 242.095000 152.760000 243.345000 ;
        RECT 150.960000 250.235000 152.760000 251.485000 ;
        RECT 129.360000 258.375000 131.160000 259.625000 ;
        RECT 118.560000 258.375000 120.360000 259.625000 ;
        RECT 118.560000 266.515000 120.360000 267.765000 ;
        RECT 129.360000 266.515000 131.160000 267.765000 ;
        RECT 150.960000 266.515000 152.760000 267.765000 ;
        RECT 150.960000 258.375000 152.760000 259.625000 ;
        RECT 140.160000 266.515000 141.960000 267.765000 ;
        RECT 140.160000 258.375000 141.960000 259.625000 ;
        RECT 107.760000 290.935000 109.560000 292.185000 ;
        RECT 96.960000 290.935000 98.760000 292.185000 ;
        RECT 86.160000 290.935000 87.960000 292.185000 ;
        RECT 96.960000 282.795000 98.760000 284.045000 ;
        RECT 96.960000 274.655000 98.760000 275.905000 ;
        RECT 86.160000 274.655000 87.960000 275.905000 ;
        RECT 86.160000 282.795000 87.960000 284.045000 ;
        RECT 107.760000 274.655000 109.560000 275.905000 ;
        RECT 107.760000 282.795000 109.560000 284.045000 ;
        RECT 96.960000 299.075000 98.760000 299.865000 ;
        RECT 86.160000 299.075000 87.960000 299.865000 ;
        RECT 107.760000 299.075000 109.560000 299.865000 ;
        RECT 150.960000 290.935000 152.760000 292.185000 ;
        RECT 140.160000 290.935000 141.960000 292.185000 ;
        RECT 129.360000 290.935000 131.160000 292.185000 ;
        RECT 118.560000 290.935000 120.360000 292.185000 ;
        RECT 118.560000 274.655000 120.360000 275.905000 ;
        RECT 118.560000 282.795000 120.360000 284.045000 ;
        RECT 129.360000 274.655000 131.160000 275.905000 ;
        RECT 129.360000 282.795000 131.160000 284.045000 ;
        RECT 140.160000 274.655000 141.960000 275.905000 ;
        RECT 140.160000 282.795000 141.960000 284.045000 ;
        RECT 150.960000 274.655000 152.760000 275.905000 ;
        RECT 150.960000 282.795000 152.760000 284.045000 ;
        RECT 118.560000 299.075000 120.360000 299.865000 ;
        RECT 129.360000 299.075000 131.160000 299.865000 ;
        RECT 140.160000 299.075000 141.960000 299.865000 ;
        RECT 150.960000 299.075000 152.760000 299.865000 ;
        RECT 194.160000 193.255000 195.960000 194.505000 ;
        RECT 194.160000 185.115000 195.960000 186.365000 ;
        RECT 194.160000 176.975000 195.960000 178.225000 ;
        RECT 194.160000 168.835000 195.960000 170.085000 ;
        RECT 194.160000 160.695000 195.960000 161.945000 ;
        RECT 172.560000 168.835000 174.360000 170.085000 ;
        RECT 161.760000 160.695000 163.560000 161.945000 ;
        RECT 161.760000 168.835000 163.560000 170.085000 ;
        RECT 172.560000 160.695000 174.360000 161.945000 ;
        RECT 183.360000 168.835000 185.160000 170.085000 ;
        RECT 183.360000 160.695000 185.160000 161.945000 ;
        RECT 161.760000 176.975000 163.560000 178.225000 ;
        RECT 161.760000 185.115000 163.560000 186.365000 ;
        RECT 161.760000 193.255000 163.560000 194.505000 ;
        RECT 172.560000 176.975000 174.360000 178.225000 ;
        RECT 172.560000 185.115000 174.360000 186.365000 ;
        RECT 172.560000 193.255000 174.360000 194.505000 ;
        RECT 183.360000 176.975000 185.160000 178.225000 ;
        RECT 183.360000 185.115000 185.160000 186.365000 ;
        RECT 183.360000 193.255000 185.160000 194.505000 ;
        RECT 204.960000 168.835000 206.760000 170.085000 ;
        RECT 204.960000 160.695000 206.760000 161.945000 ;
        RECT 215.760000 160.695000 217.560000 161.945000 ;
        RECT 226.560000 160.695000 228.360000 161.945000 ;
        RECT 215.760000 168.835000 217.560000 170.085000 ;
        RECT 226.560000 168.835000 228.360000 170.085000 ;
        RECT 204.960000 176.975000 206.760000 178.225000 ;
        RECT 204.960000 185.115000 206.760000 186.365000 ;
        RECT 204.960000 193.255000 206.760000 194.505000 ;
        RECT 215.760000 176.975000 217.560000 178.225000 ;
        RECT 226.560000 176.975000 228.360000 178.225000 ;
        RECT 215.760000 193.255000 217.560000 194.505000 ;
        RECT 215.760000 185.115000 217.560000 186.365000 ;
        RECT 226.560000 185.115000 228.360000 186.365000 ;
        RECT 226.560000 193.255000 228.360000 194.505000 ;
        RECT 194.160000 225.815000 195.960000 227.065000 ;
        RECT 194.160000 217.675000 195.960000 218.925000 ;
        RECT 194.160000 209.535000 195.960000 210.785000 ;
        RECT 194.160000 201.395000 195.960000 202.645000 ;
        RECT 161.760000 201.395000 163.560000 202.645000 ;
        RECT 161.760000 209.535000 163.560000 210.785000 ;
        RECT 172.560000 201.395000 174.360000 202.645000 ;
        RECT 172.560000 209.535000 174.360000 210.785000 ;
        RECT 183.360000 201.395000 185.160000 202.645000 ;
        RECT 183.360000 209.535000 185.160000 210.785000 ;
        RECT 161.760000 217.675000 163.560000 218.925000 ;
        RECT 161.760000 225.815000 163.560000 227.065000 ;
        RECT 172.560000 217.675000 174.360000 218.925000 ;
        RECT 172.560000 225.815000 174.360000 227.065000 ;
        RECT 183.360000 217.675000 185.160000 218.925000 ;
        RECT 183.360000 225.815000 185.160000 227.065000 ;
        RECT 204.960000 201.395000 206.760000 202.645000 ;
        RECT 204.960000 209.535000 206.760000 210.785000 ;
        RECT 215.760000 201.395000 217.560000 202.645000 ;
        RECT 215.760000 209.535000 217.560000 210.785000 ;
        RECT 226.560000 201.395000 228.360000 202.645000 ;
        RECT 226.560000 209.535000 228.360000 210.785000 ;
        RECT 204.960000 217.675000 206.760000 218.925000 ;
        RECT 204.960000 225.815000 206.760000 227.065000 ;
        RECT 215.760000 217.675000 217.560000 218.925000 ;
        RECT 215.760000 225.815000 217.560000 227.065000 ;
        RECT 226.560000 217.675000 228.360000 218.925000 ;
        RECT 226.560000 225.815000 228.360000 227.065000 ;
        RECT 248.160000 168.835000 249.960000 170.085000 ;
        RECT 237.360000 160.695000 239.160000 161.945000 ;
        RECT 237.360000 168.835000 239.160000 170.085000 ;
        RECT 248.160000 160.695000 249.960000 161.945000 ;
        RECT 269.760000 168.835000 271.560000 170.085000 ;
        RECT 269.760000 160.695000 271.560000 161.945000 ;
        RECT 258.960000 168.835000 260.760000 170.085000 ;
        RECT 258.960000 160.695000 260.760000 161.945000 ;
        RECT 237.360000 176.975000 239.160000 178.225000 ;
        RECT 237.360000 185.115000 239.160000 186.365000 ;
        RECT 237.360000 193.255000 239.160000 194.505000 ;
        RECT 248.160000 176.975000 249.960000 178.225000 ;
        RECT 248.160000 185.115000 249.960000 186.365000 ;
        RECT 248.160000 193.255000 249.960000 194.505000 ;
        RECT 258.960000 176.975000 260.760000 178.225000 ;
        RECT 258.960000 185.115000 260.760000 186.365000 ;
        RECT 258.960000 193.255000 260.760000 194.505000 ;
        RECT 269.760000 176.975000 271.560000 178.225000 ;
        RECT 269.760000 185.115000 271.560000 186.365000 ;
        RECT 269.760000 193.255000 271.560000 194.505000 ;
        RECT 291.360000 168.835000 293.160000 170.085000 ;
        RECT 291.360000 160.695000 293.160000 161.945000 ;
        RECT 280.560000 168.835000 282.360000 170.085000 ;
        RECT 280.560000 160.695000 282.360000 161.945000 ;
        RECT 301.680000 168.835000 303.680000 170.085000 ;
        RECT 301.680000 160.695000 303.680000 161.945000 ;
        RECT 291.360000 193.255000 293.160000 194.505000 ;
        RECT 291.360000 185.115000 293.160000 186.365000 ;
        RECT 291.360000 176.975000 293.160000 178.225000 ;
        RECT 280.560000 193.255000 282.360000 194.505000 ;
        RECT 280.560000 185.115000 282.360000 186.365000 ;
        RECT 280.560000 176.975000 282.360000 178.225000 ;
        RECT 301.680000 193.255000 303.680000 194.505000 ;
        RECT 301.680000 185.115000 303.680000 186.365000 ;
        RECT 301.680000 176.975000 303.680000 178.225000 ;
        RECT 237.360000 201.395000 239.160000 202.645000 ;
        RECT 237.360000 209.535000 239.160000 210.785000 ;
        RECT 248.160000 201.395000 249.960000 202.645000 ;
        RECT 248.160000 209.535000 249.960000 210.785000 ;
        RECT 258.960000 201.395000 260.760000 202.645000 ;
        RECT 258.960000 209.535000 260.760000 210.785000 ;
        RECT 269.760000 201.395000 271.560000 202.645000 ;
        RECT 269.760000 209.535000 271.560000 210.785000 ;
        RECT 237.360000 217.675000 239.160000 218.925000 ;
        RECT 237.360000 225.815000 239.160000 227.065000 ;
        RECT 248.160000 217.675000 249.960000 218.925000 ;
        RECT 248.160000 225.815000 249.960000 227.065000 ;
        RECT 258.960000 217.675000 260.760000 218.925000 ;
        RECT 258.960000 225.815000 260.760000 227.065000 ;
        RECT 269.760000 217.675000 271.560000 218.925000 ;
        RECT 269.760000 225.815000 271.560000 227.065000 ;
        RECT 291.360000 209.535000 293.160000 210.785000 ;
        RECT 291.360000 201.395000 293.160000 202.645000 ;
        RECT 280.560000 209.535000 282.360000 210.785000 ;
        RECT 280.560000 201.395000 282.360000 202.645000 ;
        RECT 301.680000 201.395000 303.680000 202.645000 ;
        RECT 301.680000 209.535000 303.680000 210.785000 ;
        RECT 291.360000 225.815000 293.160000 227.065000 ;
        RECT 291.360000 217.675000 293.160000 218.925000 ;
        RECT 280.560000 225.815000 282.360000 227.065000 ;
        RECT 280.560000 217.675000 282.360000 218.925000 ;
        RECT 301.680000 217.675000 303.680000 218.925000 ;
        RECT 301.680000 225.815000 303.680000 227.065000 ;
        RECT 194.160000 266.515000 195.960000 267.765000 ;
        RECT 194.160000 258.375000 195.960000 259.625000 ;
        RECT 194.160000 250.235000 195.960000 251.485000 ;
        RECT 194.160000 242.095000 195.960000 243.345000 ;
        RECT 194.160000 233.955000 195.960000 235.205000 ;
        RECT 161.760000 233.955000 163.560000 235.205000 ;
        RECT 161.760000 242.095000 163.560000 243.345000 ;
        RECT 161.760000 250.235000 163.560000 251.485000 ;
        RECT 172.560000 233.955000 174.360000 235.205000 ;
        RECT 172.560000 242.095000 174.360000 243.345000 ;
        RECT 172.560000 250.235000 174.360000 251.485000 ;
        RECT 183.360000 233.955000 185.160000 235.205000 ;
        RECT 183.360000 242.095000 185.160000 243.345000 ;
        RECT 183.360000 250.235000 185.160000 251.485000 ;
        RECT 172.560000 266.515000 174.360000 267.765000 ;
        RECT 161.760000 258.375000 163.560000 259.625000 ;
        RECT 161.760000 266.515000 163.560000 267.765000 ;
        RECT 172.560000 258.375000 174.360000 259.625000 ;
        RECT 183.360000 266.515000 185.160000 267.765000 ;
        RECT 183.360000 258.375000 185.160000 259.625000 ;
        RECT 204.960000 233.955000 206.760000 235.205000 ;
        RECT 204.960000 242.095000 206.760000 243.345000 ;
        RECT 204.960000 250.235000 206.760000 251.485000 ;
        RECT 215.760000 242.095000 217.560000 243.345000 ;
        RECT 215.760000 233.955000 217.560000 235.205000 ;
        RECT 226.560000 233.955000 228.360000 235.205000 ;
        RECT 226.560000 242.095000 228.360000 243.345000 ;
        RECT 215.760000 250.235000 217.560000 251.485000 ;
        RECT 226.560000 250.235000 228.360000 251.485000 ;
        RECT 204.960000 266.515000 206.760000 267.765000 ;
        RECT 204.960000 258.375000 206.760000 259.625000 ;
        RECT 215.760000 258.375000 217.560000 259.625000 ;
        RECT 226.560000 258.375000 228.360000 259.625000 ;
        RECT 215.760000 266.515000 217.560000 267.765000 ;
        RECT 226.560000 266.515000 228.360000 267.765000 ;
        RECT 194.160000 299.075000 195.960000 299.865000 ;
        RECT 194.160000 290.935000 195.960000 292.185000 ;
        RECT 194.160000 282.795000 195.960000 284.045000 ;
        RECT 194.160000 274.655000 195.960000 275.905000 ;
        RECT 183.360000 290.935000 185.160000 292.185000 ;
        RECT 172.560000 290.935000 174.360000 292.185000 ;
        RECT 161.760000 290.935000 163.560000 292.185000 ;
        RECT 161.760000 274.655000 163.560000 275.905000 ;
        RECT 161.760000 282.795000 163.560000 284.045000 ;
        RECT 172.560000 274.655000 174.360000 275.905000 ;
        RECT 172.560000 282.795000 174.360000 284.045000 ;
        RECT 183.360000 274.655000 185.160000 275.905000 ;
        RECT 183.360000 282.795000 185.160000 284.045000 ;
        RECT 183.360000 299.075000 185.160000 299.865000 ;
        RECT 172.560000 299.075000 174.360000 299.865000 ;
        RECT 161.760000 299.075000 163.560000 299.865000 ;
        RECT 226.560000 290.935000 228.360000 292.185000 ;
        RECT 215.760000 290.935000 217.560000 292.185000 ;
        RECT 204.960000 290.935000 206.760000 292.185000 ;
        RECT 204.960000 274.655000 206.760000 275.905000 ;
        RECT 204.960000 282.795000 206.760000 284.045000 ;
        RECT 215.760000 274.655000 217.560000 275.905000 ;
        RECT 215.760000 282.795000 217.560000 284.045000 ;
        RECT 226.560000 274.655000 228.360000 275.905000 ;
        RECT 226.560000 282.795000 228.360000 284.045000 ;
        RECT 204.960000 299.075000 206.760000 299.865000 ;
        RECT 215.760000 299.075000 217.560000 299.865000 ;
        RECT 226.560000 299.075000 228.360000 299.865000 ;
        RECT 237.360000 233.955000 239.160000 235.205000 ;
        RECT 237.360000 242.095000 239.160000 243.345000 ;
        RECT 237.360000 250.235000 239.160000 251.485000 ;
        RECT 248.160000 233.955000 249.960000 235.205000 ;
        RECT 248.160000 242.095000 249.960000 243.345000 ;
        RECT 248.160000 250.235000 249.960000 251.485000 ;
        RECT 258.960000 233.955000 260.760000 235.205000 ;
        RECT 258.960000 242.095000 260.760000 243.345000 ;
        RECT 258.960000 250.235000 260.760000 251.485000 ;
        RECT 269.760000 233.955000 271.560000 235.205000 ;
        RECT 269.760000 242.095000 271.560000 243.345000 ;
        RECT 269.760000 250.235000 271.560000 251.485000 ;
        RECT 248.160000 266.515000 249.960000 267.765000 ;
        RECT 237.360000 258.375000 239.160000 259.625000 ;
        RECT 237.360000 266.515000 239.160000 267.765000 ;
        RECT 248.160000 258.375000 249.960000 259.625000 ;
        RECT 269.760000 266.515000 271.560000 267.765000 ;
        RECT 269.760000 258.375000 271.560000 259.625000 ;
        RECT 258.960000 266.515000 260.760000 267.765000 ;
        RECT 258.960000 258.375000 260.760000 259.625000 ;
        RECT 291.360000 250.235000 293.160000 251.485000 ;
        RECT 291.360000 242.095000 293.160000 243.345000 ;
        RECT 291.360000 233.955000 293.160000 235.205000 ;
        RECT 280.560000 250.235000 282.360000 251.485000 ;
        RECT 280.560000 242.095000 282.360000 243.345000 ;
        RECT 280.560000 233.955000 282.360000 235.205000 ;
        RECT 301.680000 250.235000 303.680000 251.485000 ;
        RECT 301.680000 242.095000 303.680000 243.345000 ;
        RECT 301.680000 233.955000 303.680000 235.205000 ;
        RECT 291.360000 266.515000 293.160000 267.765000 ;
        RECT 291.360000 258.375000 293.160000 259.625000 ;
        RECT 280.560000 266.515000 282.360000 267.765000 ;
        RECT 280.560000 258.375000 282.360000 259.625000 ;
        RECT 301.680000 266.515000 303.680000 267.765000 ;
        RECT 301.680000 258.375000 303.680000 259.625000 ;
        RECT 269.760000 290.935000 271.560000 292.185000 ;
        RECT 258.960000 290.935000 260.760000 292.185000 ;
        RECT 248.160000 290.935000 249.960000 292.185000 ;
        RECT 237.360000 290.935000 239.160000 292.185000 ;
        RECT 237.360000 274.655000 239.160000 275.905000 ;
        RECT 237.360000 282.795000 239.160000 284.045000 ;
        RECT 248.160000 274.655000 249.960000 275.905000 ;
        RECT 248.160000 282.795000 249.960000 284.045000 ;
        RECT 258.960000 274.655000 260.760000 275.905000 ;
        RECT 258.960000 282.795000 260.760000 284.045000 ;
        RECT 269.760000 274.655000 271.560000 275.905000 ;
        RECT 269.760000 282.795000 271.560000 284.045000 ;
        RECT 237.360000 299.075000 239.160000 299.865000 ;
        RECT 248.160000 299.075000 249.960000 299.865000 ;
        RECT 258.960000 299.075000 260.760000 299.865000 ;
        RECT 269.760000 299.075000 271.560000 299.865000 ;
        RECT 291.360000 290.935000 293.160000 292.185000 ;
        RECT 280.560000 290.935000 282.360000 292.185000 ;
        RECT 301.680000 290.935000 303.680000 292.185000 ;
        RECT 291.360000 282.795000 293.160000 284.045000 ;
        RECT 291.360000 274.655000 293.160000 275.905000 ;
        RECT 280.560000 282.795000 282.360000 284.045000 ;
        RECT 280.560000 274.655000 282.360000 275.905000 ;
        RECT 301.680000 274.655000 303.680000 275.905000 ;
        RECT 301.680000 282.795000 303.680000 284.045000 ;
        RECT 291.360000 299.075000 293.160000 299.865000 ;
        RECT 280.560000 299.075000 282.360000 299.865000 ;
        RECT 300.865000 299.075000 301.245000 299.445000 ;
        RECT 301.680000 299.535000 303.680000 299.865000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 311.040000 311.540000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 311.040000 311.540000 ;
    LAYER met2 ;
      RECT 0.000000 0.000000 311.040000 311.540000 ;
    LAYER met3 ;
      RECT 0.000000 0.000000 311.040000 311.540000 ;
  END
END ldo

END LIBRARY
